magic
tech scmos
timestamp 1701512323
<< nwell >>
rect -48 8 34 35
rect 41 5 66 21
<< ntransistor >>
rect 52 -12 54 -8
rect -35 -66 -32 -49
rect -14 -66 -11 -49
rect 8 -66 11 -49
<< ptransistor >>
rect -36 15 -33 27
rect -14 15 -11 27
rect 6 15 9 27
rect 52 11 54 15
<< ndiffusion >>
rect 51 -12 52 -8
rect 54 -12 55 -8
rect -43 -57 -41 -49
rect -36 -57 -35 -49
rect -43 -66 -35 -57
rect -32 -66 -14 -49
rect -11 -66 8 -49
rect 11 -58 20 -49
rect 11 -66 26 -58
<< pdiffusion >>
rect -42 18 -41 27
rect -37 18 -36 27
rect -42 15 -36 18
rect -33 18 -27 27
rect -23 18 -14 27
rect -33 15 -14 18
rect -11 18 -5 27
rect -1 18 6 27
rect -11 15 6 18
rect 9 18 14 27
rect 18 18 26 27
rect 9 15 26 18
rect 51 11 52 15
rect 54 11 55 15
<< ndcontact >>
rect 47 -12 51 -8
rect 55 -12 59 -8
rect -41 -57 -36 -49
rect 20 -58 26 -49
<< pdcontact >>
rect -41 18 -37 27
rect -27 18 -23 27
rect -5 18 -1 27
rect 14 18 18 27
rect 47 11 51 15
rect 55 11 59 15
<< polysilicon >>
rect -36 27 -33 37
rect -14 27 -11 38
rect 6 27 9 37
rect 52 15 54 18
rect -36 3 -33 15
rect -46 0 -33 3
rect -14 -8 -11 15
rect 6 -8 9 15
rect 52 0 54 11
rect 43 -3 54 0
rect 52 -8 54 -3
rect 52 -15 54 -12
rect -35 -49 -32 -37
rect -14 -49 -11 -29
rect 8 -49 11 -29
rect -35 -70 -32 -66
rect -14 -70 -11 -66
rect 8 -70 11 -66
<< polycontact >>
rect -50 0 -46 4
rect 39 -3 43 1
rect -14 -12 -10 -8
rect 5 -12 9 -8
rect -14 -29 -10 -25
rect 8 -29 12 -25
rect -35 -37 -31 -33
<< metal1 >>
rect -41 41 53 46
rect -41 27 -37 41
rect -5 27 -1 41
rect 48 24 53 41
rect 41 21 66 24
rect -60 0 -50 4
rect -27 1 -23 18
rect 14 1 18 18
rect 47 15 51 21
rect 55 1 59 11
rect -60 -33 -56 0
rect -27 -3 39 1
rect 55 -2 82 1
rect -26 -12 -14 -8
rect -5 -12 5 -8
rect -26 -25 -21 -12
rect -5 -25 0 -12
rect -26 -29 -14 -25
rect -5 -29 8 -25
rect -60 -37 -35 -33
rect 20 -49 26 -3
rect 55 -8 59 -2
rect 47 -16 51 -12
rect 41 -21 60 -16
rect -41 -91 -36 -57
rect 48 -91 54 -21
rect -41 -95 54 -91
<< end >>
