magic
tech scmos
timestamp 1701523680
<< nwell >>
rect -3 -38 51 -11
rect 86 -41 111 -25
rect -8 -196 46 -169
rect 81 -199 106 -183
rect -11 -356 43 -329
rect 78 -359 103 -343
rect -17 -690 37 -663
rect 72 -693 97 -677
rect -22 -848 32 -821
rect 67 -851 92 -835
rect -25 -1008 29 -981
rect 64 -1011 89 -995
rect -24 -1167 30 -1140
rect 65 -1170 90 -1154
<< ntransistor >>
rect 97 -58 99 -54
rect 10 -112 13 -95
rect 23 -112 26 -95
rect 92 -216 94 -212
rect 5 -270 8 -253
rect 18 -270 21 -253
rect 89 -376 91 -372
rect 2 -430 5 -413
rect 15 -430 18 -413
rect 83 -710 85 -706
rect -4 -764 -1 -747
rect 9 -764 12 -747
rect 78 -868 80 -864
rect -9 -922 -6 -905
rect 4 -922 7 -905
rect 75 -1028 77 -1024
rect -12 -1082 -9 -1065
rect 1 -1082 4 -1065
rect 76 -1187 78 -1183
rect -11 -1241 -8 -1224
rect 2 -1241 5 -1224
<< ptransistor >>
rect 9 -31 12 -19
rect 23 -31 26 -19
rect 97 -35 99 -31
rect 4 -189 7 -177
rect 18 -189 21 -177
rect 92 -193 94 -189
rect 1 -349 4 -337
rect 15 -349 18 -337
rect 89 -353 91 -349
rect -5 -683 -2 -671
rect 9 -683 12 -671
rect 83 -687 85 -683
rect -10 -841 -7 -829
rect 4 -841 7 -829
rect 78 -845 80 -841
rect -13 -1001 -10 -989
rect 1 -1001 4 -989
rect 75 -1005 77 -1001
rect -12 -1160 -9 -1148
rect 2 -1160 5 -1148
rect 76 -1164 78 -1160
<< ndiffusion >>
rect 96 -58 97 -54
rect 99 -58 100 -54
rect 2 -103 4 -95
rect 9 -103 10 -95
rect 2 -112 10 -103
rect 13 -112 23 -95
rect 26 -103 33 -95
rect 38 -103 40 -95
rect 26 -112 40 -103
rect 91 -216 92 -212
rect 94 -216 95 -212
rect -3 -261 -1 -253
rect 4 -261 5 -253
rect -3 -270 5 -261
rect 8 -270 18 -253
rect 21 -261 28 -253
rect 33 -261 35 -253
rect 21 -270 35 -261
rect 88 -376 89 -372
rect 91 -376 92 -372
rect -6 -421 -4 -413
rect 1 -421 2 -413
rect -6 -430 2 -421
rect 5 -430 15 -413
rect 18 -421 25 -413
rect 30 -421 32 -413
rect 18 -430 32 -421
rect 82 -710 83 -706
rect 85 -710 86 -706
rect -12 -755 -10 -747
rect -5 -755 -4 -747
rect -12 -764 -4 -755
rect -1 -764 9 -747
rect 12 -755 19 -747
rect 24 -755 26 -747
rect 12 -764 26 -755
rect 77 -868 78 -864
rect 80 -868 81 -864
rect -17 -913 -15 -905
rect -10 -913 -9 -905
rect -17 -922 -9 -913
rect -6 -922 4 -905
rect 7 -913 14 -905
rect 19 -913 21 -905
rect 7 -922 21 -913
rect 74 -1028 75 -1024
rect 77 -1028 78 -1024
rect -20 -1073 -18 -1065
rect -13 -1073 -12 -1065
rect -20 -1082 -12 -1073
rect -9 -1082 1 -1065
rect 4 -1073 11 -1065
rect 16 -1073 18 -1065
rect 4 -1082 18 -1073
rect 75 -1187 76 -1183
rect 78 -1187 79 -1183
rect -19 -1232 -17 -1224
rect -12 -1232 -11 -1224
rect -19 -1241 -11 -1232
rect -8 -1241 2 -1224
rect 5 -1232 12 -1224
rect 17 -1232 19 -1224
rect 5 -1241 19 -1232
<< pdiffusion >>
rect 3 -28 4 -19
rect 8 -28 9 -19
rect 3 -31 9 -28
rect 12 -28 15 -19
rect 19 -28 23 -19
rect 12 -31 23 -28
rect 26 -28 29 -19
rect 33 -28 36 -19
rect 26 -31 36 -28
rect 96 -35 97 -31
rect 99 -35 100 -31
rect -2 -186 -1 -177
rect 3 -186 4 -177
rect -2 -189 4 -186
rect 7 -186 10 -177
rect 14 -186 18 -177
rect 7 -189 18 -186
rect 21 -186 24 -177
rect 28 -186 31 -177
rect 21 -189 31 -186
rect 91 -193 92 -189
rect 94 -193 95 -189
rect -5 -346 -4 -337
rect 0 -346 1 -337
rect -5 -349 1 -346
rect 4 -346 7 -337
rect 11 -346 15 -337
rect 4 -349 15 -346
rect 18 -346 21 -337
rect 25 -346 28 -337
rect 18 -349 28 -346
rect 88 -353 89 -349
rect 91 -353 92 -349
rect -11 -680 -10 -671
rect -6 -680 -5 -671
rect -11 -683 -5 -680
rect -2 -680 1 -671
rect 5 -680 9 -671
rect -2 -683 9 -680
rect 12 -680 15 -671
rect 19 -680 22 -671
rect 12 -683 22 -680
rect 82 -687 83 -683
rect 85 -687 86 -683
rect -16 -838 -15 -829
rect -11 -838 -10 -829
rect -16 -841 -10 -838
rect -7 -838 -4 -829
rect 0 -838 4 -829
rect -7 -841 4 -838
rect 7 -838 10 -829
rect 14 -838 17 -829
rect 7 -841 17 -838
rect 77 -845 78 -841
rect 80 -845 81 -841
rect -19 -998 -18 -989
rect -14 -998 -13 -989
rect -19 -1001 -13 -998
rect -10 -998 -7 -989
rect -3 -998 1 -989
rect -10 -1001 1 -998
rect 4 -998 7 -989
rect 11 -998 14 -989
rect 4 -1001 14 -998
rect 74 -1005 75 -1001
rect 77 -1005 78 -1001
rect -18 -1157 -17 -1148
rect -13 -1157 -12 -1148
rect -18 -1160 -12 -1157
rect -9 -1157 -6 -1148
rect -2 -1157 2 -1148
rect -9 -1160 2 -1157
rect 5 -1157 8 -1148
rect 12 -1157 15 -1148
rect 5 -1160 15 -1157
rect 75 -1164 76 -1160
rect 78 -1164 79 -1160
<< ndcontact >>
rect 92 -58 96 -54
rect 100 -58 104 -54
rect 4 -103 9 -95
rect 33 -103 38 -95
rect 87 -216 91 -212
rect 95 -216 99 -212
rect -1 -261 4 -253
rect 28 -261 33 -253
rect 84 -376 88 -372
rect 92 -376 96 -372
rect -4 -421 1 -413
rect 25 -421 30 -413
rect 78 -710 82 -706
rect 86 -710 90 -706
rect -10 -755 -5 -747
rect 19 -755 24 -747
rect 73 -868 77 -864
rect 81 -868 85 -864
rect -15 -913 -10 -905
rect 14 -913 19 -905
rect 70 -1028 74 -1024
rect 78 -1028 82 -1024
rect -18 -1073 -13 -1065
rect 11 -1073 16 -1065
rect 71 -1187 75 -1183
rect 79 -1187 83 -1183
rect -17 -1232 -12 -1224
rect 12 -1232 17 -1224
<< pdcontact >>
rect 4 -28 8 -19
rect 15 -28 19 -19
rect 29 -28 33 -19
rect 92 -35 96 -31
rect 100 -35 104 -31
rect -1 -186 3 -177
rect 10 -186 14 -177
rect 24 -186 28 -177
rect 87 -193 91 -189
rect 95 -193 99 -189
rect -4 -346 0 -337
rect 7 -346 11 -337
rect 21 -346 25 -337
rect 84 -353 88 -349
rect 92 -353 96 -349
rect -10 -680 -6 -671
rect 1 -680 5 -671
rect 15 -680 19 -671
rect 78 -687 82 -683
rect 86 -687 90 -683
rect -15 -838 -11 -829
rect -4 -838 0 -829
rect 10 -838 14 -829
rect 73 -845 77 -841
rect 81 -845 85 -841
rect -18 -998 -14 -989
rect -7 -998 -3 -989
rect 7 -998 11 -989
rect 70 -1005 74 -1001
rect 78 -1005 82 -1001
rect -17 -1157 -13 -1148
rect -6 -1157 -2 -1148
rect 8 -1157 12 -1148
rect 71 -1164 75 -1160
rect 79 -1164 83 -1160
<< polysilicon >>
rect 9 -19 12 -9
rect 23 -19 26 -8
rect 97 -31 99 -28
rect 9 -43 12 -31
rect -1 -46 12 -43
rect 23 -64 26 -31
rect 97 -46 99 -35
rect 88 -49 99 -46
rect 97 -54 99 -49
rect 97 -61 99 -58
rect 10 -95 13 -83
rect 23 -95 26 -68
rect 10 -116 13 -112
rect 23 -116 26 -112
rect 4 -177 7 -167
rect 18 -177 21 -166
rect 92 -189 94 -186
rect 4 -201 7 -189
rect -6 -204 7 -201
rect 18 -222 21 -189
rect 92 -204 94 -193
rect 83 -207 94 -204
rect 92 -212 94 -207
rect 92 -219 94 -216
rect 5 -253 8 -241
rect 18 -253 21 -226
rect 5 -274 8 -270
rect 18 -274 21 -270
rect 1 -337 4 -327
rect 15 -337 18 -326
rect 89 -349 91 -346
rect 1 -361 4 -349
rect -9 -364 4 -361
rect 15 -382 18 -349
rect 89 -364 91 -353
rect 80 -367 91 -364
rect 89 -372 91 -367
rect 89 -379 91 -376
rect 2 -413 5 -401
rect 15 -413 18 -386
rect 2 -434 5 -430
rect 15 -434 18 -430
rect -5 -671 -2 -661
rect 9 -671 12 -660
rect 83 -683 85 -680
rect -5 -695 -2 -683
rect -15 -698 -2 -695
rect 9 -716 12 -683
rect 83 -698 85 -687
rect 74 -701 85 -698
rect 83 -706 85 -701
rect 83 -713 85 -710
rect -4 -747 -1 -735
rect 9 -747 12 -720
rect -4 -768 -1 -764
rect 9 -768 12 -764
rect -10 -829 -7 -819
rect 4 -829 7 -818
rect 78 -841 80 -838
rect -10 -853 -7 -841
rect -20 -856 -7 -853
rect 4 -874 7 -841
rect 78 -856 80 -845
rect 69 -859 80 -856
rect 78 -864 80 -859
rect 78 -871 80 -868
rect -9 -905 -6 -893
rect 4 -905 7 -878
rect -9 -926 -6 -922
rect 4 -926 7 -922
rect -13 -989 -10 -979
rect 1 -989 4 -978
rect 75 -1001 77 -998
rect -13 -1013 -10 -1001
rect -23 -1016 -10 -1013
rect 1 -1034 4 -1001
rect 75 -1016 77 -1005
rect 66 -1019 77 -1016
rect 75 -1024 77 -1019
rect 75 -1031 77 -1028
rect -12 -1065 -9 -1053
rect 1 -1065 4 -1038
rect -12 -1086 -9 -1082
rect 1 -1086 4 -1082
rect -12 -1148 -9 -1138
rect 2 -1148 5 -1137
rect 76 -1160 78 -1157
rect -12 -1172 -9 -1160
rect -22 -1175 -9 -1172
rect 2 -1193 5 -1160
rect 76 -1175 78 -1164
rect 67 -1178 78 -1175
rect 76 -1183 78 -1178
rect 76 -1190 78 -1187
rect -11 -1224 -8 -1212
rect 2 -1224 5 -1197
rect -11 -1245 -8 -1241
rect 2 -1245 5 -1241
<< polycontact >>
rect -5 -46 -1 -42
rect 84 -49 88 -45
rect 23 -68 27 -64
rect 10 -83 14 -79
rect -10 -204 -6 -200
rect 79 -207 83 -203
rect 18 -226 22 -222
rect 5 -241 9 -237
rect -13 -364 -9 -360
rect 76 -367 80 -363
rect 15 -386 19 -382
rect 2 -401 6 -397
rect -19 -698 -15 -694
rect 70 -701 74 -697
rect 9 -720 13 -716
rect -4 -735 0 -731
rect -24 -856 -20 -852
rect 65 -859 69 -855
rect 4 -878 8 -874
rect -9 -893 -5 -889
rect -27 -1016 -23 -1012
rect 62 -1019 66 -1015
rect 1 -1038 5 -1034
rect -12 -1053 -8 -1049
rect -26 -1175 -22 -1171
rect 63 -1178 67 -1174
rect 2 -1197 6 -1193
rect -11 -1212 -7 -1208
<< metal1 >>
rect 51 153 58 165
rect 126 108 142 111
rect 53 7 60 18
rect 4 -5 66 0
rect 72 -5 98 0
rect 4 -19 8 -5
rect 29 -19 33 -5
rect 93 -22 98 -5
rect 86 -25 111 -22
rect -15 -46 -5 -42
rect 15 -45 19 -28
rect 92 -31 96 -25
rect 100 -45 104 -35
rect -15 -47 -11 -46
rect 15 -49 84 -45
rect 100 -48 134 -45
rect -15 -79 -11 -55
rect 20 -68 23 -64
rect -15 -83 10 -79
rect 33 -95 38 -49
rect 100 -54 104 -48
rect 4 -137 9 -103
rect 92 -137 96 -58
rect 4 -142 39 -137
rect 45 -142 96 -137
rect -1 -163 65 -158
rect 71 -163 93 -158
rect -1 -177 3 -163
rect 24 -177 28 -163
rect 88 -180 93 -163
rect 81 -183 106 -180
rect -20 -204 -10 -200
rect 10 -203 14 -186
rect 87 -189 91 -183
rect 95 -203 99 -193
rect -20 -205 -16 -204
rect 10 -207 79 -203
rect 95 -206 130 -203
rect -20 -237 -16 -213
rect 15 -226 18 -222
rect -20 -241 5 -237
rect 28 -253 33 -207
rect 95 -212 99 -206
rect -1 -295 4 -261
rect 87 -295 91 -216
rect -1 -300 41 -295
rect 47 -300 91 -295
rect -4 -323 67 -318
rect 73 -323 90 -318
rect -4 -337 0 -323
rect 21 -337 25 -323
rect 85 -340 90 -323
rect 78 -343 103 -340
rect -23 -364 -13 -360
rect 7 -363 11 -346
rect 84 -349 88 -343
rect 92 -363 96 -353
rect -23 -365 -19 -364
rect 7 -367 76 -363
rect 92 -366 128 -363
rect -23 -397 -19 -373
rect 12 -386 15 -382
rect -23 -401 2 -397
rect 25 -413 30 -367
rect 92 -372 96 -366
rect -4 -455 1 -421
rect 84 -455 88 -376
rect -4 -460 38 -455
rect 44 -460 88 -455
rect -10 -657 65 -652
rect 71 -657 84 -652
rect -10 -671 -6 -657
rect 15 -671 19 -657
rect 79 -674 84 -657
rect 72 -677 97 -674
rect -29 -698 -19 -694
rect 1 -697 5 -680
rect 78 -683 82 -677
rect 86 -697 90 -687
rect -29 -699 -25 -698
rect 1 -701 70 -697
rect 86 -700 121 -697
rect -29 -731 -25 -707
rect 6 -720 9 -716
rect -29 -735 -4 -731
rect 19 -747 24 -701
rect 86 -706 90 -700
rect -10 -789 -5 -755
rect 78 -789 82 -710
rect -10 -794 39 -789
rect 45 -794 82 -789
rect -15 -815 65 -810
rect 71 -815 79 -810
rect -15 -829 -11 -815
rect 10 -829 14 -815
rect 74 -832 79 -815
rect 67 -835 92 -832
rect -34 -856 -24 -852
rect -4 -855 0 -838
rect 73 -841 77 -835
rect 81 -855 85 -845
rect -34 -857 -30 -856
rect -4 -859 65 -855
rect 81 -858 118 -855
rect -34 -889 -30 -865
rect 1 -878 4 -874
rect -34 -893 -9 -889
rect 14 -905 19 -859
rect 81 -864 85 -858
rect -15 -947 -10 -913
rect 73 -947 77 -868
rect -15 -952 40 -947
rect 46 -952 77 -947
rect -18 -975 65 -970
rect -18 -989 -14 -975
rect 7 -989 11 -975
rect 71 -992 76 -970
rect 64 -995 89 -992
rect -37 -1016 -27 -1012
rect -7 -1015 -3 -998
rect 70 -1001 74 -995
rect 78 -1015 82 -1005
rect -37 -1017 -33 -1016
rect -7 -1019 62 -1015
rect 78 -1018 116 -1015
rect -37 -1049 -33 -1025
rect -2 -1038 1 -1034
rect -37 -1053 -12 -1049
rect 11 -1065 16 -1019
rect 78 -1024 82 -1018
rect -18 -1107 -13 -1073
rect 70 -1107 74 -1028
rect -18 -1112 39 -1107
rect 45 -1112 74 -1107
rect -17 -1134 65 -1129
rect 71 -1134 77 -1129
rect -17 -1148 -13 -1134
rect 8 -1148 12 -1134
rect 72 -1151 77 -1134
rect 65 -1154 90 -1151
rect -36 -1175 -26 -1171
rect -6 -1174 -2 -1157
rect 71 -1160 75 -1154
rect 79 -1174 83 -1164
rect -36 -1176 -32 -1175
rect -6 -1178 63 -1174
rect 79 -1177 114 -1174
rect -36 -1208 -32 -1184
rect -1 -1197 2 -1193
rect -36 -1212 -11 -1208
rect 12 -1224 17 -1178
rect 79 -1183 83 -1177
rect -17 -1266 -12 -1232
rect 71 -1266 75 -1187
rect -17 -1271 39 -1266
rect 45 -1271 75 -1266
<< m2contact >>
rect 66 151 72 156
rect -14 96 -6 104
rect 16 82 25 92
rect 37 14 43 19
rect 66 -5 72 0
rect -19 -55 -11 -47
rect 11 -73 20 -64
rect 39 -142 45 -137
rect 65 -163 71 -158
rect -24 -213 -16 -205
rect 6 -231 15 -222
rect 41 -300 47 -295
rect 67 -323 73 -318
rect -27 -373 -19 -365
rect 3 -391 12 -382
rect 38 -460 44 -455
rect 65 -657 71 -652
rect -33 -707 -25 -699
rect -3 -725 6 -716
rect 39 -794 45 -789
rect 65 -815 71 -810
rect -38 -865 -30 -857
rect -8 -883 1 -874
rect 40 -952 46 -947
rect 65 -975 71 -970
rect -41 -1025 -33 -1017
rect -11 -1043 -2 -1034
rect 39 -1112 45 -1107
rect 65 -1134 71 -1129
rect -40 -1184 -32 -1176
rect -10 -1202 -1 -1193
rect 39 -1271 45 -1266
<< metal2 >>
rect -175 92 -165 152
rect -89 96 -14 104
rect -175 82 16 92
rect -175 -63 -165 82
rect 37 19 49 169
rect 43 14 49 19
rect -97 -55 -19 -47
rect -175 -64 -96 -63
rect -175 -73 11 -64
rect 20 -73 23 -64
rect -175 -83 -165 -73
rect -175 -221 -164 -83
rect 37 -137 49 14
rect 37 -142 39 -137
rect 45 -142 49 -137
rect -102 -213 -24 -205
rect -175 -222 -99 -221
rect -175 -231 6 -222
rect 15 -231 18 -222
rect -175 -382 -164 -231
rect 37 -295 49 -142
rect 37 -300 41 -295
rect 47 -300 49 -295
rect -105 -373 -27 -365
rect -175 -391 3 -382
rect 12 -391 15 -382
rect -175 -392 -99 -391
rect -175 -716 -164 -392
rect 37 -455 49 -300
rect 37 -460 38 -455
rect 44 -460 49 -455
rect -111 -707 -33 -699
rect -175 -725 -3 -716
rect 6 -725 9 -716
rect -175 -726 -100 -725
rect -175 -807 -164 -726
rect -176 -873 -164 -807
rect 37 -789 49 -460
rect 37 -794 39 -789
rect 45 -794 49 -789
rect -116 -865 -38 -857
rect -176 -874 -101 -873
rect -176 -883 -8 -874
rect 1 -883 4 -874
rect -176 -891 -164 -883
rect -176 -1035 -165 -891
rect 37 -947 49 -794
rect 37 -952 40 -947
rect 46 -952 49 -947
rect -119 -1025 -41 -1017
rect -120 -1035 -11 -1034
rect -176 -1043 -11 -1035
rect -2 -1043 1 -1034
rect -176 -1045 -101 -1043
rect -176 -1193 -165 -1045
rect 37 -1107 49 -952
rect 37 -1112 39 -1107
rect 45 -1112 49 -1107
rect -118 -1184 -40 -1176
rect -176 -1202 -10 -1193
rect -1 -1202 2 -1193
rect -176 -1212 -165 -1202
rect 37 -1266 49 -1112
rect 37 -1271 39 -1266
rect 45 -1271 49 -1266
rect 37 -1277 49 -1271
rect 63 156 75 169
rect 63 151 66 156
rect 72 151 75 156
rect 63 0 75 151
rect 63 -5 66 0
rect 72 -5 75 0
rect 63 -158 75 -5
rect 63 -163 65 -158
rect 71 -163 75 -158
rect 63 -318 75 -163
rect 63 -323 67 -318
rect 73 -323 75 -318
rect 63 -652 75 -323
rect 63 -657 65 -652
rect 71 -657 75 -652
rect 63 -810 75 -657
rect 63 -815 65 -810
rect 71 -815 75 -810
rect 63 -970 75 -815
rect 63 -975 65 -970
rect 71 -975 75 -970
rect 63 -1129 75 -975
rect 63 -1134 65 -1129
rect 71 -1134 75 -1129
rect 63 -1277 75 -1134
use AND  AND_0
timestamp 1700315882
transform 1 0 50 0 1 110
box -60 -96 78 46
<< labels >>
rlabel metal1 109 -1177 112 -1174 1 b3_out
rlabel metal1 109 -1018 112 -1015 1 b2_out
rlabel metal1 110 -858 113 -855 1 b1_out
rlabel metal1 111 -700 114 -697 1 b0_out
rlabel metal1 121 -366 124 -363 1 a3_out
rlabel metal1 123 -206 126 -203 1 a2_out
rlabel metal1 125 -48 128 -45 1 a1_out
rlabel metal1 139 108 142 111 7 a0_out
<< end >>
