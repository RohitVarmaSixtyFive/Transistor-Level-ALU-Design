* SPICE3 file created from not.ext - technology: scmos

.option scale=0.09u
.include TSMC_180nm.txt
.global gnd
.param SUPPLY = 1.8

Vdd VDD gnd 'SUPPLY'

V_in_a A gnd PULSE(0 1.8 0ns 100ps 100ps 50ns 70ns)

M1000 out A VDD w_n9_1# CMOSP w=4 l=2
+  ad=20 pd=18 as=20 ps=18
M1001 out A gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=20 ps=18
C0 out gnd 0.08fF
C1 VDD out 0.07fF
C2 VDD w_n9_1# 0.05fF
C3 out A 0.02fF
C4 w_n9_1# A 0.06fF
C5 gnd A 0.01fF
C6 out w_n9_1# 0.03fF
C7 gnd Gnd 0.08fF
C8 out Gnd 0.06fF
C9 VDD Gnd 0.04fF
C10 A Gnd 0.17fF
C11 w_n9_1# Gnd 0.40fF

.tran 1n 1000n
.measure tran trise0 
+ TRIG v(A) VAL = 'SUPPLY/2' RISE =1
+ TARG v(out) VAL = 'SUPPLY/2' FALL =1 

.measure tran tfall0
+ TRIG v(A) VAL = 'SUPPLY/2' FALL =1 
+ TARG v(out) VAL = 'SUPPLY/2' RISE=1

.measure tran tpd_A param = '(trise0 + tfall0)/2' goal = 0
* .measure tran trise1
* + TRIG v(w2) VAL = 'SUPPLout/2' RISE =1
* + TARG v(out) VAL = 'SUPPLout/2' FALL =1 

* .measure tran tfall1
* + TRIG v(w2) VAL = 'SUPPLout/2' FALL =1 
* + TARG v(out) VAL = 'SUPPLout/2' RISE=1

* .measure tran tpd_w2 param = '(trise1 + tfall1)/2' goal = 0
.control
run
plot v(A) v(out)+2
* hardcopy image.ps v(A)
.end
.endc
