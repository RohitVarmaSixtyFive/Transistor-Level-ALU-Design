magic
tech scmos
timestamp 1701527625
<< metal1 >>
rect -35 189 -29 190
rect -35 184 99 189
rect 105 187 112 206
rect -35 55 -29 184
rect 211 141 237 144
rect -9 118 78 123
rect -77 33 -55 37
rect -9 36 -5 118
rect -33 33 -5 36
rect -77 32 -59 33
rect -72 -16 -54 -12
rect -34 -16 -29 -13
rect -72 -84 -60 -16
rect -73 -162 -60 -84
rect -31 -93 -27 -28
rect -9 -154 -5 33
rect 209 -8 235 -5
rect -9 -159 79 -154
rect 210 -158 236 -155
rect -74 -175 -59 -162
rect -74 -184 -28 -175
rect -50 -349 -40 -184
rect 206 -318 232 -315
rect -50 -359 -40 -358
rect 122 -424 126 -410
<< m2contact >>
rect 175 184 183 190
rect -53 55 -48 60
rect 104 118 111 125
rect -85 31 -77 37
rect 148 47 156 54
rect -42 16 -37 21
rect -53 6 -48 11
rect -29 -16 -24 -11
rect -42 -32 -37 -27
rect -31 -98 -25 -93
rect 175 15 183 21
rect 73 -29 78 -24
rect 101 -30 107 -24
rect 90 -98 98 -91
rect 148 -101 156 -94
rect 175 -135 181 -130
rect -28 -184 -15 -172
rect 102 -184 112 -174
rect 148 -252 156 -245
rect 175 -275 181 -269
rect 69 -336 78 -327
rect 99 -342 108 -334
rect -50 -358 -40 -349
rect 148 -412 156 -405
<< metal2 >>
rect 9 118 104 125
rect -85 -33 -78 31
rect -53 11 -49 55
rect -42 -27 -38 16
rect 9 -11 14 118
rect -31 -16 -29 -11
rect -24 -16 14 -11
rect 8 -24 14 -16
rect 8 -29 73 -24
rect 101 -33 107 -30
rect -85 -35 -74 -33
rect -86 -43 -74 -35
rect 5 -39 107 -33
rect 5 -43 13 -39
rect -86 -49 13 -43
rect -86 -327 -74 -49
rect -25 -98 90 -93
rect 148 -94 156 47
rect 175 21 181 184
rect 175 14 181 15
rect -15 -183 102 -174
rect 112 -183 118 -174
rect 148 -245 156 -101
rect 176 -130 181 14
rect -86 -336 69 -327
rect 78 -336 79 -327
rect 99 -349 108 -342
rect -40 -358 108 -349
rect 148 -405 156 -252
rect 175 -269 181 -135
rect 175 -290 181 -275
use NOT  NOT_0
timestamp 1700315584
transform 1 0 -47 0 1 -11
box -9 -20 16 20
use NOT  NOT_1
timestamp 1700315584
transform 1 0 -48 0 1 38
box -9 -20 16 20
use AND  AND_0
timestamp 1700315882
transform 1 0 135 0 1 143
box -60 -96 78 46
use AND  AND_1
timestamp 1700315882
transform 1 0 134 0 1 -6
box -60 -96 78 46
use AND  AND_2
timestamp 1700315882
transform 1 0 136 0 1 -156
box -60 -96 78 46
use AND  AND_3
timestamp 1700315882
transform 1 0 134 0 1 -316
box -60 -96 78 46
<< labels >>
rlabel metal1 224 -318 228 -315 1 d3
rlabel metal1 220 -158 224 -155 1 d2
rlabel metal1 217 -8 221 -5 1 d1
rlabel metal1 223 141 227 144 1 d0
<< end >>
