* SPICE3 file created from four_or.ext - technology: scmos
.include TSMC_180nm.txt

.param SUPPLY = 1.8

.global gnd

Vdd VDD gnd 'SUPPLY'

V_in_a a gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)
V_in_b b gnd PULSE(1.8 0 0ns 100ps 100ps 100ns 100ns)
V_in_c c gnd PULSE(1.8 0 0ns 100ps 100ps 100ns 200s)
V_in_d d gnd PULSE(1.8 0 0ns 100ps 100ps 100ns 300ns)

.option scale=0.09u

M1000 gnd c in Gnd CMOSN w=4 l=2
+  ad=116 pd=78 as=88 ps=68
M1001 in d a_7_9# VDD CMOSP w=4 l=2
+  ad=20 pd=18 as=32 ps=24
M1002 in b gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 out in gnd Gnd CMOSN w=6 l=2
+  ad=42 pd=26 as=0 ps=0
M1004 in d gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 a_n5_9# b a_n16_9# VDD CMOSP w=4 l=2
+  ad=40 pd=28 as=36 ps=26
M1006 out in VDD VDD CMOSP w=6 l=2
+  ad=42 pd=26 as=68 ps=46
M1007 a_7_9# c a_n5_9# VDD CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 a_n16_9# a VDD VDD CMOSP w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1009 gnd a in Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
C0 out gnd 0.05fF
C1 in b 0.06fF
C2 VDD VDD 0.09fF
C3 gnd c 0.05fF
C4 in VDD 0.09fF
C5 c b 0.01fF
C6 out VDD 0.03fF
C7 VDD a 0.06fF
C8 VDD VDD 0.09fF
C9 in a 0.06fF
C10 VDD d 0.07fF
C11 gnd b 0.04fF
C12 in d 0.26fF
C13 VDD in 0.04fF
C14 out in 0.07fF
C15 VDD in 0.07fF
C16 VDD c 0.07fF
C17 VDD out 0.03fF
C18 gnd a 0.05fF
C19 in c 0.06fF
C20 gnd d 0.04fF
C21 in gnd 0.33fF
C22 VDD b 0.07fF
C23 gnd Gnd 0.41fF
C24 out Gnd 0.16fF
C25 VDD Gnd 0.21fF
C26 in Gnd 0.37fF
C27 d Gnd 0.33fF
C28 c Gnd 0.27fF
C29 b Gnd 0.26fF
C30 a Gnd 0.31fF
C31 VDD Gnd 1.02fF
C32 VDD Gnd 1.07fF
.tran 1n 1000n

* .measure tran trise0 
* + TRIG v(A) VAL = 'SUPPLY/2' FALL =1
* + TARG v(OUT) VAL = 'SUPPLY/2' RISE =1 

* .measure tran tfall0
* + TRIG v(A) VAL = 'SUPPLY/2' RISE =1 
* + TARG v(OUT) VAL = 'SUPPLY/2' FALL=1

* .measure tran tpd_a_b0 param = '(trise0 + tfall0)/2' goal = 0

.control
run
* set color0 = rgb:f/f/e
* set color1 = white
plot v(a) v(b)+2 v(c)+4 v(d)+6 v(out)+8
* plot v(OUT_FINAL)/
* hardcopy image.ps v(node_a) v(node_b)+2 v(node_out)+4
.end
.endc