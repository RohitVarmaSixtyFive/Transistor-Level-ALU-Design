magic
tech scmos
timestamp 1699296593
<< nwell >>
rect -48 8 63 35
rect 130 5 155 21
<< ntransistor >>
rect 141 -12 143 -8
rect -35 -66 -32 -49
rect -14 -66 -11 -49
rect 8 -66 11 -49
rect 32 -66 35 -49
rect 54 -66 57 -49
<< ptransistor >>
rect -36 15 -33 27
rect -14 15 -11 27
rect 6 15 9 27
rect 26 15 29 27
rect 46 15 49 27
rect 141 11 143 15
<< ndiffusion >>
rect 140 -12 141 -8
rect 143 -12 144 -8
rect -43 -57 -41 -49
rect -36 -57 -35 -49
rect -43 -66 -35 -57
rect -32 -66 -14 -49
rect -11 -66 8 -49
rect 11 -66 32 -49
rect 35 -66 54 -49
rect 57 -57 59 -49
rect 64 -57 65 -49
rect 57 -66 65 -57
<< pdiffusion >>
rect -42 18 -41 27
rect -37 18 -36 27
rect -42 15 -36 18
rect -33 18 -27 27
rect -23 18 -14 27
rect -33 15 -14 18
rect -11 18 -5 27
rect -1 18 6 27
rect -11 15 6 18
rect 9 18 14 27
rect 18 18 26 27
rect 9 15 26 18
rect 29 18 38 27
rect 42 18 46 27
rect 29 15 46 18
rect 49 18 50 27
rect 54 18 57 27
rect 49 15 57 18
rect 140 11 141 15
rect 143 11 144 15
<< ndcontact >>
rect 136 -12 140 -8
rect 144 -12 148 -8
rect -41 -57 -36 -49
rect 59 -57 64 -49
<< pdcontact >>
rect -41 18 -37 27
rect -27 18 -23 27
rect -5 18 -1 27
rect 14 18 18 27
rect 38 18 42 27
rect 50 18 54 27
rect 136 11 140 15
rect 144 11 148 15
<< polysilicon >>
rect -36 27 -33 37
rect -14 27 -11 38
rect 6 27 9 37
rect 26 27 29 38
rect 46 27 49 38
rect 141 15 143 18
rect -36 3 -33 15
rect -46 0 -33 3
rect -14 -8 -11 15
rect 6 -8 9 15
rect 26 -8 29 15
rect 46 6 49 15
rect 46 3 56 6
rect 52 -8 56 3
rect 141 0 143 11
rect 132 -3 143 0
rect 141 -8 143 -3
rect 141 -15 143 -12
rect 56 -28 57 -24
rect -35 -49 -32 -37
rect -14 -49 -11 -29
rect 8 -49 11 -29
rect 32 -49 35 -29
rect 54 -49 57 -28
rect -35 -70 -32 -66
rect -14 -70 -11 -66
rect 8 -70 11 -66
rect 32 -70 35 -66
rect 54 -70 57 -66
<< polycontact >>
rect -50 0 -46 4
rect -14 -12 -10 -8
rect 5 -12 9 -8
rect 128 -3 132 1
rect 26 -12 30 -8
rect 52 -12 56 -8
rect -14 -29 -10 -25
rect 8 -29 12 -25
rect 31 -29 35 -25
rect 52 -28 56 -24
rect -35 -37 -31 -33
<< metal1 >>
rect -41 41 142 46
rect -41 27 -37 41
rect -5 27 -1 41
rect 38 27 42 41
rect 137 24 142 41
rect 130 21 155 24
rect -60 0 -50 4
rect -27 2 -23 18
rect 14 2 18 18
rect 50 2 54 18
rect 136 15 140 21
rect -27 1 132 2
rect -60 -33 -56 0
rect -27 -2 128 1
rect -26 -12 -14 -8
rect -5 -12 5 -8
rect 19 -12 26 -8
rect 39 -12 52 -8
rect -26 -25 -21 -12
rect -5 -25 0 -12
rect 19 -25 24 -12
rect 39 -24 44 -12
rect -26 -29 -14 -25
rect -5 -29 8 -25
rect 19 -29 31 -25
rect 39 -28 52 -24
rect -60 -37 -35 -33
rect 59 -49 64 -2
rect 144 1 148 11
rect 144 -2 162 1
rect 144 -8 148 -2
rect 136 -16 140 -12
rect 130 -21 149 -16
rect -41 -91 -36 -57
rect 137 -91 143 -21
rect -41 -99 151 -91
<< labels >>
rlabel metal1 -58 0 -56 4 3 a
rlabel metal1 -26 -21 -21 -16 1 b
rlabel metal1 -5 -20 0 -15 1 c
rlabel metal1 19 -22 24 -17 1 d
rlabel metal1 39 -21 44 -16 1 e
rlabel metal1 152 -2 155 1 1 out
rlabel polycontact 128 -3 132 1 1 in
rlabel metal1 83 -97 89 -93 1 gnd
rlabel metal1 105 43 106 44 5 VDD
<< end >>
