magic
tech scmos
timestamp 1701545641
<< polysilicon >>
rect 553 591 558 2973
rect 909 2906 1421 2920
rect 797 1556 832 1563
rect 797 1360 804 1556
rect 855 1388 859 1418
rect 855 1387 986 1388
rect 1654 1387 1658 1417
rect 855 1384 2273 1387
rect 982 1383 2273 1384
rect 797 1353 917 1360
rect 910 1236 917 1353
rect 982 1159 986 1383
rect 962 1155 986 1159
rect 2269 1046 2273 1383
rect 2269 1042 2449 1046
rect 868 556 873 610
rect 264 551 873 556
rect 386 409 390 470
rect 263 405 390 409
rect 2960 378 2990 382
rect 2960 345 2964 378
rect 2736 341 2964 345
rect 315 -1955 319 281
rect 2736 -5 2740 341
rect 2736 -9 2982 -5
rect 814 -63 841 -56
rect 814 -285 821 -63
rect 875 -263 879 -201
rect 875 -267 996 -263
rect 814 -292 931 -285
rect 924 -402 931 -292
rect 992 -475 996 -267
rect 970 -476 996 -475
rect 975 -479 996 -476
rect 2978 -619 2982 -9
rect 2391 -623 2982 -619
rect 1208 -906 1234 -895
rect 1208 -959 1219 -906
rect 1042 -970 1219 -959
rect 1208 -1100 1224 -1071
rect 1043 -1101 1224 -1100
rect 1055 -1116 1224 -1101
rect 1066 -1214 1214 -1213
rect 1075 -1222 1214 -1214
rect 2391 -1955 2395 -623
rect 315 -1959 2395 -1955
<< polycontact >>
rect 553 2973 566 2983
rect 894 2906 909 2923
rect 832 1555 840 1563
rect 855 1418 860 1423
rect 1654 1417 1659 1422
rect 910 1226 918 1236
rect 956 1153 962 1159
rect 868 610 873 615
rect 553 583 561 591
rect 259 551 264 556
rect 386 470 391 476
rect 258 405 263 410
rect 2990 378 2996 383
rect 841 -64 849 -56
rect 875 -201 880 -196
rect 924 -409 931 -402
rect 970 -481 975 -476
rect 1234 -906 1245 -895
rect 1031 -970 1042 -959
rect 1208 -1071 1224 -1058
rect 1043 -1116 1055 -1101
rect 1066 -1222 1075 -1214
rect 1214 -1222 1220 -1209
<< metal1 >>
rect 553 2983 1172 2984
rect 566 2973 1172 2983
rect 894 2885 908 2906
rect 182 2878 908 2885
rect 182 641 189 2878
rect 901 2847 908 2878
rect 1161 2807 1172 2973
rect 989 2797 1138 2800
rect 445 1628 671 1637
rect 173 635 189 641
rect 182 634 189 635
rect 260 606 381 611
rect 310 508 314 579
rect 374 528 381 606
rect 310 504 353 508
rect 446 501 450 1628
rect 743 707 754 2315
rect 759 1177 764 2785
rect 1135 2770 1138 2797
rect 1161 2796 1271 2807
rect 1296 2791 1299 2849
rect 1288 2788 1299 2791
rect 1288 2770 1291 2788
rect 1135 2767 1291 2770
rect 1029 2734 1254 2740
rect 774 2642 781 2643
rect 742 694 754 696
rect 311 497 366 501
rect 431 497 450 501
rect 168 482 174 487
rect -15 466 -6 472
rect 311 433 317 497
rect 553 433 559 583
rect 311 427 560 433
rect -14 418 7 423
rect 315 280 319 281
rect 310 277 684 280
rect 299 -456 302 120
rect 299 -459 698 -456
rect 742 -932 747 694
rect 759 -463 764 1166
rect 774 1023 781 2634
rect 774 -614 781 1015
rect 789 865 796 2484
rect 1029 1992 1032 2734
rect 968 1989 1032 1992
rect 1057 1834 1060 2650
rect 961 1831 1060 1834
rect 1094 1674 1097 2576
rect 956 1671 1097 1674
rect 1141 1515 1144 2516
rect 960 1512 1144 1515
rect 2213 1478 2410 1482
rect 2406 1197 2410 1478
rect 990 1178 1910 1181
rect 988 1022 1819 1025
rect 983 864 1738 867
rect 789 856 796 857
rect 791 -772 794 856
rect 981 704 1689 707
rect 1686 222 1689 704
rect 1735 333 1738 864
rect 1816 407 1819 1022
rect 1907 487 1910 1178
rect 1955 407 1958 642
rect 1816 404 1958 407
rect 1987 333 1990 565
rect 3098 398 3107 401
rect 2942 389 2966 392
rect 2942 369 2945 389
rect 2714 366 2945 369
rect 1735 330 1990 333
rect 1685 217 1689 222
rect 1685 213 2051 217
rect 1264 -425 1283 -423
rect 971 -430 1283 -425
rect 1264 -431 1283 -430
rect 1000 -459 1165 -456
rect 970 -476 975 -475
rect 993 -615 1135 -612
rect 998 -773 1110 -770
rect 995 -933 1090 -930
rect 1032 -1264 1035 -970
rect 987 -1267 1035 -1264
rect 1043 -1422 1046 -1116
rect 984 -1425 1046 -1422
rect 1067 -1582 1070 -1222
rect 1087 -1346 1090 -933
rect 1107 -1197 1110 -773
rect 1132 -1042 1135 -615
rect 1162 -880 1165 -459
rect 1275 -834 1283 -431
rect 1365 -879 1373 -876
rect 1162 -883 1220 -880
rect 1365 -1027 1381 -1024
rect 1132 -1045 1208 -1042
rect 1362 -1178 1377 -1175
rect 1107 -1198 1206 -1197
rect 1107 -1200 1210 -1198
rect 1363 -1329 1372 -1326
rect 1087 -1349 1202 -1346
rect 1208 -1349 1209 -1346
rect 983 -1585 1070 -1582
rect 1174 -1361 1218 -1358
rect 1174 -1741 1177 -1361
rect 983 -1744 1177 -1741
rect 1256 -1833 1261 -1418
rect 929 -1838 1261 -1833
<< m2contact >>
rect 759 2785 767 2793
rect 742 2315 754 2324
rect 671 1623 686 1637
rect 1271 2796 1282 2807
rect 1254 2734 1262 2741
rect 774 2634 782 2642
rect 979 2641 984 2646
rect 757 1166 767 1177
rect 742 696 754 707
rect 684 275 696 286
rect 698 -459 708 -450
rect 774 1015 782 1023
rect 758 -471 766 -463
rect 976 2483 981 2488
rect 975 2323 980 2328
rect 1057 2650 1067 2660
rect 1093 2576 1103 2586
rect 1140 2516 1150 2526
rect 1259 2441 1267 2450
rect 1249 2066 1259 2075
rect 1308 1655 1315 1662
rect 789 857 797 865
rect 774 -622 781 -614
rect 976 370 982 376
rect 1954 642 1962 651
rect 2076 642 2084 651
rect 1907 479 1915 487
rect 1987 565 1993 571
rect 2063 565 2069 571
rect 2088 479 2095 486
rect 972 212 979 219
rect 971 52 978 59
rect 969 -107 976 -100
rect 791 -780 800 -772
rect 740 -940 748 -932
rect 1208 -1047 1213 -1042
rect 1246 -1047 1251 -1042
rect 1206 -1198 1212 -1192
rect 1243 -1198 1249 -1192
rect 1202 -1349 1208 -1343
rect 1244 -1349 1250 -1343
<< metal2 >>
rect 2053 2837 2061 2841
rect 1270 2796 1271 2807
rect 732 2785 759 2793
rect 767 2785 770 2793
rect 1067 2657 1261 2660
rect 733 2634 758 2642
rect 984 2641 991 2646
rect 986 2510 991 2641
rect 1103 2578 1262 2581
rect 1150 2520 1219 2523
rect 986 2505 1173 2510
rect 729 2476 755 2484
rect 981 2483 1000 2488
rect 995 2358 1000 2483
rect 1168 2446 1173 2505
rect 1216 2504 1219 2520
rect 1216 2501 1260 2504
rect 1168 2441 1259 2446
rect 1267 2441 1269 2446
rect 2051 2441 2064 2445
rect 1168 2438 1173 2441
rect 995 2353 1256 2358
rect 720 2316 742 2324
rect 754 2316 758 2324
rect 980 2323 1024 2328
rect 1018 2006 1023 2323
rect 1251 2075 1256 2353
rect 2047 2045 2067 2050
rect 1018 2001 1313 2006
rect 724 1982 741 1990
rect 720 1824 739 1832
rect 717 1664 736 1672
rect 1308 1662 1313 2001
rect 2041 1619 2070 1623
rect 722 1506 741 1514
rect 2233 1455 2246 1459
rect 767 1166 773 1174
rect 1962 642 2076 651
rect 1993 565 2063 571
rect 1915 479 2088 486
rect 1058 471 2041 474
rect 1058 377 1061 471
rect 975 376 1061 377
rect 975 374 976 376
rect 982 374 1061 376
rect 1348 368 2020 372
rect 1348 238 1352 368
rect 974 234 1352 238
rect 1476 283 2018 286
rect 974 219 978 234
rect 1476 75 1479 283
rect 2015 281 2018 283
rect 976 72 1479 75
rect 1602 202 2027 205
rect 976 59 979 72
rect 978 52 979 59
rect 968 -105 969 -102
rect 1602 -102 1605 202
rect 976 -105 1605 -102
rect 744 -471 758 -463
rect 766 -471 789 -463
rect 748 -940 781 -932
rect 1213 -1047 1246 -1042
rect 1212 -1198 1243 -1192
rect 742 -1273 745 -1266
rect 754 -1273 780 -1266
rect 754 -1274 772 -1273
rect 1208 -1349 1244 -1343
<< m3contact >>
rect 745 1981 754 1990
rect 758 1824 767 1832
rect 778 1663 787 1671
rect 799 1504 808 1512
rect 745 363 754 372
rect 758 205 767 213
rect 778 45 787 53
rect 799 -114 808 -106
rect 745 -1273 754 -1266
rect 758 -1432 767 -1423
rect 778 -1592 787 -1583
rect 800 -1751 810 -1742
<< metal3 >>
rect 745 372 754 1981
rect 745 -1266 754 363
rect 758 213 767 1824
rect 758 -1423 767 205
rect 778 53 787 1663
rect 778 -1583 787 45
rect 799 1512 808 1513
rect 799 -106 808 1504
rect 799 -1273 808 -114
rect 800 -1742 807 -1273
use comparator  comparator_0
timestamp 1701545641
transform 1 0 2108 0 1 433
box -93 -926 713 768
use AND  AND_0
timestamp 1700315882
transform 1 0 3023 0 1 400
box -60 -96 78 46
use aluand  aluand_0
timestamp 1701532374
transform 1 0 1219 0 1 -979
box -7 -445 147 157
use adder_subtractor  adder_subtractor_0
timestamp 1701531472
transform 1 0 1285 0 1 2700
box -50 -1305 949 223
use 2_input_OR  2_input_OR_0
timestamp 1701467916
transform 1 0 366 0 1 494
box -23 -24 68 39
use enable_out  enable_out_2
timestamp 1701523680
transform 1 0 873 0 1 -567
box -176 -1277 142 169
use enable_out  enable_out_1
timestamp 1701523680
transform 1 0 859 0 1 1070
box -176 -1277 142 169
use enable_out  enable_out_0
timestamp 1701523680
transform 1 0 850 0 1 2689
box -176 -1277 142 169
use decoder  decoder_0
timestamp 1701527625
transform 1 0 77 0 1 435
box -86 -424 237 206
<< labels >>
rlabel metal2 735 2787 738 2790 1 a0
rlabel metal2 734 2636 735 2638 1 a1
rlabel metal2 732 2479 733 2481 1 a2
rlabel metal2 723 2319 725 2320 1 a3
rlabel metal2 725 1983 726 1986 1 b0
rlabel metal2 721 1826 722 1827 1 b1
rlabel metal2 718 1667 719 1668 1 b2
rlabel metal2 723 1508 724 1509 1 b3
rlabel metal1 -13 467 -11 470 3 s0
rlabel metal1 -13 420 -12 421 3 s1
rlabel metal1 175 637 178 639 1 vdd
rlabel metal1 168 483 169 485 1 gnd
rlabel metal1 1166 2796 1175 2803 1 d1_decoder_wala
rlabel metal1 3105 398 3106 400 7 equal_to
rlabel metal2 2058 2838 2059 2839 1 as0
rlabel metal2 2060 2442 2063 2444 1 as1
rlabel metal2 2059 2047 2062 2048 1 as2
rlabel metal2 2061 1620 2066 1622 1 as3
rlabel metal2 2242 1456 2244 1458 1 as_carry
rlabel metal1 1370 -878 1371 -877 1 and_out0
rlabel metal1 1374 -1026 1378 -1025 1 and_out1
rlabel metal1 1372 -1177 1375 -1176 1 and_out2
rlabel metal1 1367 -1329 1370 -1327 1 and_out3
<< end >>
