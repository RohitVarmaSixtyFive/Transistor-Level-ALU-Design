* SPICE3 file created from five_and.ext - technology: scmos

.include TSMC_180nm.txt


.param SUPPLY = 1.8


.global gnd

Vdd VDD gnd 'SUPPLY'

V_in_a a gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)
* V_in_b b gnd PULSE(0 1.8 0ns 100ps 100ps 40ns 90ns)
V_in_b b gnd DC 1.8

* V_in_c c gnd PULSE(0 1.8 0ns 100ps 100ps 40ns 80ns)
V_in_c c gnd DC 1.8
* V_in_d d gnd PULSE(0 1.8 0ns 100ps 100ps 60ns 120ns)
V_in_d d gnd DC 1.8
* V_in_e e gnd PULSE(0 1.8 0ns 100ps 100ps 70ns 140ns)
V_in_e e gnd DC 1.8

.option scale=0.09u

M1000 a_35_n66# d a_11_n66# Gnd CMOSN w=17 l=3
+  ad=323 pd=72 as=357 ps=76
M1001 VDD d in VDD CMOSP w=12 l=3
+  ad=500 pd=170 as=528 ps=160
M1002 in a VDD VDD CMOSP w=12 l=3
+  ad=0 pd=0 as=0 ps=0
M1003 out in VDD VDD CMOSP w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1004 VDD b in VDD CMOSP w=12 l=3
+  ad=0 pd=0 as=0 ps=0
M1005 a_n11_n66# b a_n32_n66# Gnd CMOSN w=17 l=3
+  ad=323 pd=72 as=306 ps=70
M1006 in e VDD VDD CMOSP w=12 l=3
+  ad=0 pd=0 as=0 ps=0
M1007 a_n32_n66# a gnd Gnd CMOSN w=17 l=3
+  ad=0 pd=0 as=156 ps=68
M1008 a_11_n66# c a_n11_n66# Gnd CMOSN w=17 l=3
+  ad=0 pd=0 as=0 ps=0
M1009 in c VDD VDD CMOSP w=12 l=3
+  ad=0 pd=0 as=0 ps=0
M1010 out in gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1011 in e a_35_n66# Gnd CMOSN w=17 l=3
+  ad=136 pd=50 as=0 ps=0
C0 VDD c 0.11fF
C1 VDD in 0.08fF
C2 e d 0.03fF
C3 d c 0.02fF
C4 VDD b 0.11fF
C5 d in 0.17fF
C6 VDD a 0.11fF
C7 VDD d 0.11fF
C8 e in 0.41fF
C9 out VDD 0.07fF
C10 c in 0.19fF
C11 VDD VDD 0.05fF
C12 VDD in 0.06fF
C13 out VDD 0.03fF
C14 c b 0.07fF
C15 b in 0.20fF
C16 gnd out 0.08fF
C17 e VDD 0.11fF
C18 VDD VDD 0.08fF
C19 gnd Gnd 1.33fF
C20 out Gnd 0.09fF
C21 in Gnd 0.88fF
C22 VDD Gnd 0.82fF
C23 e Gnd 0.60fF
C24 d Gnd 0.17fF
C25 c Gnd 0.18fF
C26 b Gnd 0.53fF
C27 a Gnd 0.12fF
C28 VDD Gnd 0.03fF
C29 VDD Gnd 3.01fF
.tran 1n 1000n

.measure tran tfall0 
+ TRIG v(a) VAL = 'SUPPLY/2' FALL =1
+ TARG v(out) VAL = 'SUPPLY/2' FALL =1 

.measure tran trise0
+ TRIG v(a) VAL = 'SUPPLY/2' RISE =1 
+ TARG v(out) VAL = 'SUPPLY/2' RISE=1

.measure tran tpd_a param = '(trise0 + tfall0)/2' goal = 0

* .measure tran trise1
* + TRIG v(b) VAL = 'SUPPLY/2' RISE =1
* + TARG v(out) VAL = 'SUPPLY/2' FALL =1 

* .measure tran tfall1
* + TRIG v(b) VAL = 'SUPPLY/2' FALL =1 
* + TARG v(out) VAL = 'SUPPLY/2' RISE=1

* .measure tran tpd_b param = '(trise1 + tfall1)/2' goal = 0

* .measure tran trise2
* + TRIG v(c) VAL = 'SUPPLY/2' RISE =1
* + TARG v(out) VAL = 'SUPPLY/2' FALL =1 

* .measure tran tfall2
* + TRIG v(c) VAL = 'SUPPLY/2' FALL =1 
* + TARG v(out) VAL = 'SUPPLY/2' RISE=1

* .measure tran tpd_c param = '(trise2 + tfall2)/2' goal = 0

* .measure tran trise3
* + TRIG v(d) VAL = 'SUPPLY/2' RISE =1
* + TARG v(out) VAL = 'SUPPLY/2' FALL =1 

* .measure tran tfall3
* + TRIG v(d) VAL = 'SUPPLY/2' FALL =1 
* + TARG v(out) VAL = 'SUPPLY/2' RISE=1

* .measure tran tpd_d param = '(trise3 + tfall3)/2' goal = 0

* .measure tran trise4
* + TRIG v(e) VAL = 'SUPPLY/2' RISE =1
* + TARG v(out) VAL = 'SUPPLY/2' FALL =1 

* .measure tran tfall4
* + TRIG v(e) VAL = 'SUPPLY/2' FALL =1 
* + TARG v(out) VAL = 'SUPPLY/2' RISE=1

* .measure tran tpd_e param = '(trise4 + tfall4)/2' goal = 0

.control
run
* set color0 = rgb:f/f/e
* set color1 = white
plot v(a) v(b)+2 v(c)+4 v(d)+6 v(e)+8 v(out)+10
* plot v(OUT_FINAL)/
* hardcopy image.ps v(node_a) v(node_b)+2 v(node_out)+4
.end
.endc