* SPICE3 file created from 3_AND.ext - technology: scmos
.include TSMC_180nm.txt

.param SUPPLY = 1.8

.global gnd

Vdd VDD gnd 'SUPPLY'

V_in_a a gnd PULSE(1.8 0 0ns 100ps 100ps 40ns 100ns)
V_in_b b gnd PULSE(1.8 0 0ns 100ps 100ps 40ns 100ns)
V_in_c c gnd PULSE(1.8 0 0ns 100ps 100ps 40ns 100ns)
V_in_d d gnd PULSE(1.8 0 0ns 100ps 100ps 40ns 100ns)

.option scale=0.01u

M1000 out a_n33_15# vdd w_94_5# CMOSP w=36 l=18
+  ad=1620 pd=162 as=39528 ps=1512
M1001 out a_n33_15# gnd Gnd CMOSN w=36 l=18
+  ad=1620 pd=162 as=12636 ps=612
M1002 a_n33_15# d a_11_n66# Gnd CMOSN w=153 l=27
+  ad=13770 pd=486 as=28917 ps=684
M1003 vdd d a_n33_15# w_n48_8# CMOSP w=108 l=27
+  ad=0 pd=0 as=34992 ps=1080
M1004 a_n33_15# a vdd w_n48_8# CMOSP w=108 l=27
+  ad=0 pd=0 as=0 ps=0
M1005 vdd b a_n33_15# w_n48_8# CMOSP w=108 l=27
+  ad=0 pd=0 as=0 ps=0
M1006 a_n11_n66# b a_n32_n66# Gnd CMOSN w=153 l=27
+  ad=26163 pd=648 as=24786 ps=630
M1007 a_n32_n66# a gnd Gnd CMOSN w=153 l=27
+  ad=0 pd=0 as=0 ps=0
M1008 a_11_n66# c a_n11_n66# Gnd CMOSN w=153 l=27
+  ad=0 pd=0 as=0 ps=0
M1009 a_n33_15# c vdd w_n48_8# CMOSP w=108 l=27
+  ad=0 pd=0 as=0 ps=0

.tran 1n 1000n

* .measure tran trise0 
* + TRIG v(A) VAL = 'SUPPLY/2' FALL =1
* + TARG v(OUT) VAL = 'SUPPLY/2' RISE =1 

* .measure tran tfall0
* + TRIG v(A) VAL = 'SUPPLY/2' RISE =1 
* + TARG v(OUT) VAL = 'SUPPLY/2' FALL=1

* .measure tran tpd_a_b0 param = '(trise0 + tfall0)/2' goal = 0

.control
run
* set color0 = rgb:f/f/e
* set color1 = white
plot v(a) v(b)+2 v(c)+4 v(d)+6 v(out)+8
* plot v(OUT_FINAL)/
* hardcopy image.ps v(node_a) v(node_b)+2 v(node_out)+4
.end
.endc