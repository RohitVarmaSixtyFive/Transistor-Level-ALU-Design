magic
tech scmos
timestamp 1701339318
<< nwell >>
rect -12 10 14 27
rect 20 10 73 27
rect 79 10 105 27
<< ntransistor >>
rect 0 -11 2 -6
rect 32 -11 34 -6
rect 40 -11 42 -6
rect 50 -11 52 -6
rect 58 -11 60 -6
rect 90 -11 92 -6
<< ptransistor >>
rect 0 16 2 21
rect 32 16 34 21
rect 40 16 42 21
rect 50 16 52 21
rect 58 16 60 21
rect 90 16 92 21
<< ndiffusion >>
rect -2 -11 0 -6
rect 2 -11 4 -6
rect 31 -11 32 -6
rect 34 -11 35 -6
rect 39 -11 40 -6
rect 42 -11 43 -6
rect 47 -11 50 -6
rect 52 -11 53 -6
rect 57 -11 58 -6
rect 60 -11 62 -6
rect 67 -11 68 -6
rect 89 -11 90 -6
rect 92 -11 93 -6
<< pdiffusion >>
rect -2 16 0 21
rect 2 16 4 21
rect 26 16 27 21
rect 31 16 32 21
rect 34 16 40 21
rect 42 16 43 21
rect 47 16 50 21
rect 52 16 58 21
rect 60 16 62 21
rect 66 16 67 21
rect 89 16 90 21
rect 92 16 93 21
rect 97 16 99 21
<< ndcontact >>
rect -6 -11 -2 -6
rect 4 -11 8 -6
rect 26 -11 31 -6
rect 35 -11 39 -6
rect 43 -11 47 -6
rect 53 -11 57 -6
rect 62 -11 67 -6
rect 85 -11 89 -6
rect 93 -11 97 -6
<< pdcontact >>
rect -6 16 -2 21
rect 4 16 8 21
rect 27 16 31 21
rect 43 16 47 21
rect 62 16 66 21
rect 85 16 89 21
rect 93 16 97 21
<< polysilicon >>
rect 15 29 52 31
rect 0 21 2 24
rect 15 20 19 29
rect 32 21 34 24
rect 40 21 42 24
rect 50 21 52 29
rect 58 29 92 31
rect 58 21 60 29
rect 90 21 92 29
rect 0 8 2 16
rect 1 4 2 8
rect 0 -6 2 4
rect 32 -6 34 16
rect 40 -6 42 16
rect 50 -6 52 16
rect 58 -6 60 16
rect 0 -13 2 -11
rect 32 -13 34 -11
rect 0 -15 34 -13
rect 40 -17 42 -11
rect 50 -14 52 -11
rect 58 -14 60 -11
rect 70 -17 72 4
rect 90 -6 92 16
rect 90 -14 92 -11
rect 40 -19 72 -17
<< polycontact >>
rect 15 16 19 20
rect -3 4 1 8
rect 69 4 73 8
rect 92 2 96 6
<< metal1 >>
rect -13 33 105 37
rect -6 21 -2 33
rect 27 21 31 33
rect 62 21 66 33
rect 93 21 97 33
rect 4 9 8 16
rect 15 9 19 16
rect -18 4 -3 8
rect 4 5 19 9
rect 43 8 47 16
rect 43 7 61 8
rect 4 -6 8 5
rect 35 4 61 7
rect 85 8 89 16
rect 73 4 89 8
rect 35 3 66 4
rect 26 -6 31 -5
rect 35 -6 39 3
rect 43 -6 47 -5
rect 62 -6 67 -5
rect 85 -6 89 4
rect 96 2 100 6
rect -6 -28 -2 -11
rect 53 -28 57 -11
rect 93 -28 97 -11
rect -13 -32 105 -28
<< m2contact >>
rect 61 4 66 9
rect 26 -5 31 0
rect 43 -5 48 0
rect 62 -5 67 0
rect 100 1 105 6
<< metal2 >>
rect 77 10 116 14
rect 77 9 82 10
rect 66 4 81 9
rect -20 -5 -9 -2
rect 31 -4 43 0
rect 48 -4 62 0
rect -13 -21 -9 -5
rect 101 -21 105 1
rect -13 -25 105 -21
<< end >>
