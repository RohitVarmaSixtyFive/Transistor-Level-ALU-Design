magic
tech scmos
timestamp 1701531472
<< nwell >>
rect 14 -28 40 -11
rect 46 -28 99 -11
rect 105 -28 131 -11
rect 15 -107 41 -90
rect 47 -107 100 -90
rect 106 -107 132 -90
rect 16 -184 42 -167
rect 48 -184 101 -167
rect 107 -184 133 -167
<< ntransistor >>
rect 26 -49 28 -44
rect 58 -49 60 -44
rect 66 -49 68 -44
rect 76 -49 78 -44
rect 84 -49 86 -44
rect 116 -49 118 -44
rect 27 -128 29 -123
rect 59 -128 61 -123
rect 67 -128 69 -123
rect 77 -128 79 -123
rect 85 -128 87 -123
rect 117 -128 119 -123
rect 28 -205 30 -200
rect 60 -205 62 -200
rect 68 -205 70 -200
rect 78 -205 80 -200
rect 86 -205 88 -200
rect 118 -205 120 -200
<< ptransistor >>
rect 26 -22 28 -17
rect 58 -22 60 -17
rect 66 -22 68 -17
rect 76 -22 78 -17
rect 84 -22 86 -17
rect 116 -22 118 -17
rect 27 -101 29 -96
rect 59 -101 61 -96
rect 67 -101 69 -96
rect 77 -101 79 -96
rect 85 -101 87 -96
rect 117 -101 119 -96
rect 28 -178 30 -173
rect 60 -178 62 -173
rect 68 -178 70 -173
rect 78 -178 80 -173
rect 86 -178 88 -173
rect 118 -178 120 -173
<< ndiffusion >>
rect 24 -49 26 -44
rect 28 -49 30 -44
rect 57 -49 58 -44
rect 60 -49 61 -44
rect 65 -49 66 -44
rect 68 -49 69 -44
rect 73 -49 76 -44
rect 78 -49 79 -44
rect 83 -49 84 -44
rect 86 -49 88 -44
rect 93 -49 94 -44
rect 115 -49 116 -44
rect 118 -49 119 -44
rect 25 -128 27 -123
rect 29 -128 31 -123
rect 58 -128 59 -123
rect 61 -128 62 -123
rect 66 -128 67 -123
rect 69 -128 70 -123
rect 74 -128 77 -123
rect 79 -128 80 -123
rect 84 -128 85 -123
rect 87 -128 89 -123
rect 94 -128 95 -123
rect 116 -128 117 -123
rect 119 -128 120 -123
rect 26 -205 28 -200
rect 30 -205 32 -200
rect 59 -205 60 -200
rect 62 -205 63 -200
rect 67 -205 68 -200
rect 70 -205 71 -200
rect 75 -205 78 -200
rect 80 -205 81 -200
rect 85 -205 86 -200
rect 88 -205 90 -200
rect 95 -205 96 -200
rect 117 -205 118 -200
rect 120 -205 121 -200
<< pdiffusion >>
rect 24 -22 26 -17
rect 28 -22 30 -17
rect 52 -22 53 -17
rect 57 -22 58 -17
rect 60 -22 66 -17
rect 68 -22 69 -17
rect 73 -22 76 -17
rect 78 -22 84 -17
rect 86 -22 88 -17
rect 92 -22 93 -17
rect 115 -22 116 -17
rect 118 -22 119 -17
rect 123 -22 125 -17
rect 25 -101 27 -96
rect 29 -101 31 -96
rect 53 -101 54 -96
rect 58 -101 59 -96
rect 61 -101 67 -96
rect 69 -101 70 -96
rect 74 -101 77 -96
rect 79 -101 85 -96
rect 87 -101 89 -96
rect 93 -101 94 -96
rect 116 -101 117 -96
rect 119 -101 120 -96
rect 124 -101 126 -96
rect 26 -178 28 -173
rect 30 -178 32 -173
rect 54 -178 55 -173
rect 59 -178 60 -173
rect 62 -178 68 -173
rect 70 -178 71 -173
rect 75 -178 78 -173
rect 80 -178 86 -173
rect 88 -178 90 -173
rect 94 -178 95 -173
rect 117 -178 118 -173
rect 120 -178 121 -173
rect 125 -178 127 -173
<< ndcontact >>
rect 20 -49 24 -44
rect 30 -49 34 -44
rect 52 -49 57 -44
rect 61 -49 65 -44
rect 69 -49 73 -44
rect 79 -49 83 -44
rect 88 -49 93 -44
rect 111 -49 115 -44
rect 119 -49 123 -44
rect 21 -128 25 -123
rect 31 -128 35 -123
rect 53 -128 58 -123
rect 62 -128 66 -123
rect 70 -128 74 -123
rect 80 -128 84 -123
rect 89 -128 94 -123
rect 112 -128 116 -123
rect 120 -128 124 -123
rect 22 -205 26 -200
rect 32 -205 36 -200
rect 54 -205 59 -200
rect 63 -205 67 -200
rect 71 -205 75 -200
rect 81 -205 85 -200
rect 90 -205 95 -200
rect 113 -205 117 -200
rect 121 -205 125 -200
<< pdcontact >>
rect 20 -22 24 -17
rect 30 -22 34 -17
rect 53 -22 57 -17
rect 69 -22 73 -17
rect 88 -22 92 -17
rect 111 -22 115 -17
rect 119 -22 123 -17
rect 21 -101 25 -96
rect 31 -101 35 -96
rect 54 -101 58 -96
rect 70 -101 74 -96
rect 89 -101 93 -96
rect 112 -101 116 -96
rect 120 -101 124 -96
rect 22 -178 26 -173
rect 32 -178 36 -173
rect 55 -178 59 -173
rect 71 -178 75 -173
rect 90 -178 94 -173
rect 113 -178 117 -173
rect 121 -178 125 -173
<< polysilicon >>
rect 128 213 387 217
rect 128 80 133 213
rect 132 76 133 80
rect 41 -9 78 -7
rect 26 -17 28 -14
rect 41 -18 45 -9
rect 58 -17 60 -14
rect 66 -17 68 -14
rect 76 -17 78 -9
rect 84 -9 118 -7
rect 84 -17 86 -9
rect 116 -17 118 -9
rect 26 -30 28 -22
rect 27 -34 28 -30
rect 26 -44 28 -34
rect 58 -44 60 -22
rect 66 -44 68 -22
rect 76 -44 78 -22
rect 84 -44 86 -22
rect 26 -51 28 -49
rect 58 -51 60 -49
rect 26 -53 60 -51
rect 66 -55 68 -49
rect 76 -52 78 -49
rect 84 -52 86 -49
rect 96 -55 98 -34
rect 116 -44 118 -22
rect 116 -52 118 -49
rect 66 -57 98 -55
rect 127 -66 131 11
rect 131 -70 176 -66
rect 42 -88 79 -86
rect 27 -96 29 -93
rect 42 -97 46 -88
rect 59 -96 61 -93
rect 67 -96 69 -93
rect 77 -96 79 -88
rect 85 -88 119 -86
rect 85 -96 87 -88
rect 117 -96 119 -88
rect 27 -109 29 -101
rect 28 -113 29 -109
rect 27 -123 29 -113
rect 59 -123 61 -101
rect 67 -123 69 -101
rect 77 -123 79 -101
rect 85 -123 87 -101
rect 27 -130 29 -128
rect 59 -130 61 -128
rect 27 -132 61 -130
rect 67 -134 69 -128
rect 77 -131 79 -128
rect 85 -131 87 -128
rect 97 -134 99 -113
rect 117 -123 119 -101
rect 117 -131 119 -128
rect 67 -136 99 -134
rect 127 -145 131 -70
rect 43 -165 80 -163
rect 28 -173 30 -170
rect 43 -174 47 -165
rect 60 -173 62 -170
rect 68 -173 70 -170
rect 78 -173 80 -165
rect 86 -165 120 -163
rect 86 -173 88 -165
rect 118 -173 120 -165
rect 28 -186 30 -178
rect 29 -190 30 -186
rect 28 -200 30 -190
rect 60 -200 62 -178
rect 68 -200 70 -178
rect 78 -200 80 -178
rect 86 -200 88 -178
rect 28 -207 30 -205
rect 60 -207 62 -205
rect 28 -209 62 -207
rect 68 -211 70 -205
rect 78 -208 80 -205
rect 86 -208 88 -205
rect 98 -211 100 -190
rect 118 -200 120 -178
rect 118 -208 120 -205
rect 68 -213 100 -211
rect 129 -222 132 -149
rect 266 -179 273 213
rect 266 -183 388 -179
rect 266 -574 273 -183
rect 570 -242 576 -60
rect 266 -578 385 -574
rect 390 -578 391 -574
rect 266 -1001 273 -578
rect 565 -637 573 -456
rect 266 -1005 380 -1001
rect 385 -1005 391 -1001
rect 562 -1066 569 -851
rect 568 -1070 569 -1066
<< polycontact >>
rect 387 213 392 217
rect 128 76 132 80
rect 127 11 131 15
rect 41 -22 45 -18
rect 23 -34 27 -30
rect 95 -34 99 -30
rect 118 -36 122 -32
rect 127 -70 131 -66
rect 176 -70 180 -66
rect 42 -101 46 -97
rect 24 -113 28 -109
rect 96 -113 100 -109
rect 119 -115 123 -111
rect 127 -149 132 -145
rect 43 -178 47 -174
rect 25 -190 29 -186
rect 97 -190 101 -186
rect 120 -192 124 -188
rect 570 -60 576 -55
rect 388 -183 393 -179
rect 129 -226 133 -222
rect 570 -248 576 -242
rect 565 -456 573 -451
rect 385 -578 390 -574
rect 565 -643 573 -637
rect 562 -851 569 -846
rect 380 -1005 385 -1001
rect 562 -1070 568 -1066
<< metal1 >>
rect -29 143 317 149
rect 69 77 73 83
rect 132 76 139 80
rect -18 47 -8 51
rect -3 47 9 51
rect -18 -30 -14 47
rect 135 -1 139 76
rect 13 -5 139 -1
rect 20 -17 24 -5
rect 53 -17 57 -5
rect 88 -17 92 -5
rect 119 -17 123 -5
rect 30 -29 34 -22
rect 41 -29 45 -22
rect -18 -34 23 -30
rect 30 -33 45 -29
rect 69 -30 73 -22
rect 69 -31 87 -30
rect -18 -109 -14 -34
rect 30 -44 34 -33
rect 61 -34 87 -31
rect 111 -30 115 -22
rect 99 -34 115 -30
rect 61 -35 92 -34
rect 52 -44 57 -43
rect 61 -44 65 -35
rect 69 -44 73 -43
rect 88 -44 93 -43
rect 111 -44 115 -34
rect 122 -36 126 -32
rect 20 -66 24 -49
rect 79 -66 83 -49
rect 119 -66 123 -49
rect 13 -70 127 -66
rect 135 -80 139 -5
rect 366 -65 375 -60
rect 176 -66 375 -65
rect 180 -70 375 -66
rect 14 -84 139 -80
rect 21 -96 25 -84
rect 54 -96 58 -84
rect 89 -96 93 -84
rect 120 -96 124 -84
rect 31 -108 35 -101
rect 42 -108 46 -101
rect -18 -113 24 -109
rect 31 -112 46 -108
rect 70 -109 74 -101
rect 70 -110 88 -109
rect -18 -186 -14 -113
rect 31 -123 35 -112
rect 62 -113 88 -110
rect 112 -109 116 -101
rect 100 -113 116 -109
rect 62 -114 93 -113
rect 53 -123 58 -122
rect 62 -123 66 -114
rect 70 -123 74 -122
rect 89 -123 94 -122
rect 112 -123 116 -113
rect 123 -115 127 -111
rect 21 -145 25 -128
rect 80 -145 84 -128
rect 120 -145 124 -128
rect 14 -149 127 -145
rect 135 -157 139 -84
rect 15 -161 139 -157
rect 22 -173 26 -161
rect 55 -173 59 -161
rect 90 -173 94 -161
rect 121 -173 125 -161
rect 32 -185 36 -178
rect 43 -185 47 -178
rect -50 -190 25 -186
rect 32 -189 47 -185
rect 71 -186 75 -178
rect 71 -187 89 -186
rect -50 -1286 -45 -190
rect 32 -200 36 -189
rect 63 -190 89 -187
rect 113 -186 117 -178
rect 101 -190 117 -186
rect 63 -191 94 -190
rect 54 -200 59 -199
rect 63 -200 67 -191
rect 71 -200 75 -199
rect 90 -200 95 -199
rect 113 -200 117 -190
rect 124 -192 128 -188
rect 22 -222 26 -205
rect 81 -222 85 -205
rect 121 -222 125 -205
rect 15 -226 129 -222
rect 70 -228 73 -226
rect -30 -259 316 -253
rect -32 -633 314 -627
rect -38 -1045 310 -1039
rect 770 -1226 817 -1219
rect 787 -1251 818 -1247
rect 787 -1256 792 -1251
rect 774 -1283 777 -1277
rect 772 -1287 816 -1283
<< m2contact >>
rect -8 47 -3 52
rect 87 -34 92 -29
rect 52 -43 57 -38
rect 69 -43 74 -38
rect 88 -43 93 -38
rect 126 -37 131 -32
rect 791 -39 797 -34
rect 88 -113 93 -108
rect 53 -122 58 -117
rect 70 -122 75 -117
rect 89 -122 94 -117
rect 127 -116 132 -111
rect 89 -190 94 -185
rect 54 -199 59 -194
rect 71 -199 76 -194
rect 90 -199 95 -194
rect 128 -193 133 -188
rect 794 -436 799 -430
rect 787 -831 796 -825
rect -50 -1291 -45 -1286
<< metal2 >>
rect 745 137 770 141
rect -9 119 301 125
rect -8 52 -3 119
rect 140 53 336 57
rect -28 38 7 41
rect 103 -28 273 -24
rect 103 -29 108 -28
rect 92 -34 107 -29
rect -28 -43 17 -40
rect 57 -42 69 -38
rect 74 -42 88 -38
rect 13 -59 17 -43
rect 127 -59 131 -37
rect 13 -63 131 -59
rect 104 -107 231 -103
rect 104 -108 109 -107
rect 93 -113 108 -108
rect -27 -122 18 -119
rect 58 -121 70 -117
rect 75 -121 89 -117
rect 14 -138 18 -122
rect 128 -138 132 -116
rect 14 -142 132 -138
rect 105 -184 211 -180
rect 105 -185 110 -184
rect 94 -190 109 -185
rect -29 -199 19 -196
rect 59 -198 71 -194
rect 76 -198 90 -194
rect 15 -215 19 -199
rect 129 -215 133 -193
rect 15 -219 133 -215
rect 206 -1135 211 -184
rect 226 -712 231 -107
rect 268 -315 273 -28
rect 791 -136 797 -39
rect 297 -142 797 -136
rect 297 -276 303 -142
rect 743 -259 768 -255
rect 268 -319 337 -315
rect 794 -538 799 -436
rect 294 -543 799 -538
rect 294 -671 301 -543
rect 740 -654 765 -650
rect 226 -717 334 -712
rect 787 -973 796 -831
rect 675 -974 816 -973
rect 290 -981 816 -974
rect 290 -1098 294 -981
rect 733 -1081 758 -1077
rect 206 -1140 330 -1135
rect 944 -1245 949 -1241
rect -50 -1300 -45 -1291
rect 806 -1300 811 -1257
rect -50 -1305 811 -1300
use XOR  XOR_1
timestamp 1701339318
transform 1 0 829 0 1 -1255
box -20 -32 116 37
use XOR  XOR_0
timestamp 1701339318
transform 1 0 26 0 1 43
box -20 -32 116 37
use full_adder  full_adder_0
timestamp 1701468074
transform 1 0 366 0 1 167
box -69 -251 429 56
use full_adder  full_adder_1
timestamp 1701468074
transform 1 0 367 0 1 -229
box -69 -251 429 56
use full_adder  full_adder_2
timestamp 1701468074
transform 1 0 363 0 1 -624
box -69 -251 429 56
use full_adder  full_adder_3
timestamp 1701468074
transform 1 0 359 0 1 -1051
box -69 -251 429 56
<< labels >>
rlabel metal1 -16 48 -14 50 3 m
rlabel metal2 -26 39 -25 40 3 b0
rlabel metal2 -25 -42 -24 -41 3 b1
rlabel metal2 -25 -121 -24 -120 3 b2
rlabel metal2 -26 -198 -25 -197 3 b3
rlabel metal1 -25 145 -22 146 1 a0
rlabel metal1 -25 -257 -22 -256 1 a1
rlabel metal1 -26 -630 -23 -629 1 a2
rlabel metal1 -30 -1044 -24 -1041 1 a3
rlabel metal2 767 138 768 139 1 s0
rlabel metal2 766 -258 767 -257 1 s1
rlabel metal2 758 -653 759 -652 1 s2
rlabel metal2 756 -1080 757 -1079 1 s3
rlabel metal2 947 -1244 948 -1242 7 carry
<< end >>
