magic
tech scmos
timestamp 1701468074
<< nwell >>
rect 228 -30 254 -13
rect 260 -30 313 -13
rect 319 -30 345 -13
rect 179 -123 233 -96
rect 268 -126 293 -110
<< ntransistor >>
rect 240 -51 242 -46
rect 272 -51 274 -46
rect 280 -51 282 -46
rect 290 -51 292 -46
rect 298 -51 300 -46
rect 330 -51 332 -46
rect 279 -143 281 -139
rect 192 -197 195 -180
rect 205 -197 208 -180
<< ptransistor >>
rect 240 -24 242 -19
rect 272 -24 274 -19
rect 280 -24 282 -19
rect 290 -24 292 -19
rect 298 -24 300 -19
rect 330 -24 332 -19
rect 191 -116 194 -104
rect 205 -116 208 -104
rect 279 -120 281 -116
<< ndiffusion >>
rect 238 -51 240 -46
rect 242 -51 244 -46
rect 271 -51 272 -46
rect 274 -51 275 -46
rect 279 -51 280 -46
rect 282 -51 283 -46
rect 287 -51 290 -46
rect 292 -51 293 -46
rect 297 -51 298 -46
rect 300 -51 302 -46
rect 307 -51 308 -46
rect 329 -51 330 -46
rect 332 -51 333 -46
rect 278 -143 279 -139
rect 281 -143 282 -139
rect 184 -188 186 -180
rect 191 -188 192 -180
rect 184 -197 192 -188
rect 195 -197 205 -180
rect 208 -188 215 -180
rect 220 -188 222 -180
rect 208 -197 222 -188
<< pdiffusion >>
rect 238 -24 240 -19
rect 242 -24 244 -19
rect 266 -24 267 -19
rect 271 -24 272 -19
rect 274 -24 280 -19
rect 282 -24 283 -19
rect 287 -24 290 -19
rect 292 -24 298 -19
rect 300 -24 302 -19
rect 306 -24 307 -19
rect 329 -24 330 -19
rect 332 -24 333 -19
rect 337 -24 339 -19
rect 185 -113 186 -104
rect 190 -113 191 -104
rect 185 -116 191 -113
rect 194 -113 197 -104
rect 201 -113 205 -104
rect 194 -116 205 -113
rect 208 -113 211 -104
rect 215 -113 218 -104
rect 208 -116 218 -113
rect 278 -120 279 -116
rect 281 -120 282 -116
<< ndcontact >>
rect 234 -51 238 -46
rect 244 -51 248 -46
rect 266 -51 271 -46
rect 275 -51 279 -46
rect 283 -51 287 -46
rect 293 -51 297 -46
rect 302 -51 307 -46
rect 325 -51 329 -46
rect 333 -51 337 -46
rect 274 -143 278 -139
rect 282 -143 286 -139
rect 186 -188 191 -180
rect 215 -188 220 -180
<< pdcontact >>
rect 234 -24 238 -19
rect 244 -24 248 -19
rect 267 -24 271 -19
rect 283 -24 287 -19
rect 302 -24 306 -19
rect 325 -24 329 -19
rect 333 -24 337 -19
rect 186 -113 190 -104
rect 197 -113 201 -104
rect 211 -113 215 -104
rect 274 -120 278 -116
rect 282 -120 286 -116
<< polysilicon >>
rect 255 -11 292 -9
rect 240 -19 242 -16
rect 255 -20 259 -11
rect 272 -19 274 -16
rect 280 -19 282 -16
rect 290 -19 292 -11
rect 298 -11 332 -9
rect 298 -19 300 -11
rect 330 -19 332 -11
rect 240 -32 242 -24
rect 241 -36 242 -32
rect 240 -46 242 -36
rect 272 -46 274 -24
rect 280 -46 282 -24
rect 290 -46 292 -24
rect 298 -46 300 -24
rect 240 -53 242 -51
rect 272 -53 274 -51
rect 240 -55 274 -53
rect 280 -57 282 -51
rect 290 -54 292 -51
rect 298 -54 300 -51
rect 310 -57 312 -36
rect 330 -46 332 -24
rect 330 -54 332 -51
rect 280 -59 312 -57
rect 191 -104 194 -94
rect 205 -104 208 -93
rect 279 -116 281 -113
rect 191 -128 194 -116
rect 181 -131 194 -128
rect 205 -149 208 -116
rect 279 -131 281 -120
rect 270 -134 281 -131
rect 279 -139 281 -134
rect 279 -146 281 -143
rect 192 -180 195 -168
rect 205 -180 208 -153
rect 192 -201 195 -197
rect 205 -201 208 -197
<< polycontact >>
rect 255 -24 259 -20
rect 237 -36 241 -32
rect 309 -36 313 -32
rect 332 -38 336 -34
rect 177 -131 181 -127
rect 266 -134 270 -130
rect 205 -153 209 -149
rect 192 -168 196 -164
<< metal1 >>
rect 87 47 93 56
rect 136 46 238 50
rect 144 23 149 27
rect 157 23 224 27
rect 9 19 20 21
rect -55 15 20 19
rect -55 -73 -49 15
rect -57 -166 -49 -73
rect -36 8 10 12
rect -36 -70 -29 8
rect 51 -63 58 -15
rect 136 -19 209 -15
rect 119 -27 128 -26
rect -36 -79 -29 -77
rect 119 -81 128 -35
rect 150 -72 193 -66
rect 203 -68 209 -19
rect 220 -32 224 23
rect 232 -3 238 46
rect 232 -7 365 -3
rect 234 -19 238 -7
rect 267 -19 271 -7
rect 302 -19 306 -7
rect 333 -19 337 -7
rect 244 -31 248 -24
rect 255 -31 259 -24
rect 220 -36 237 -32
rect 244 -35 259 -31
rect 283 -32 287 -24
rect 283 -33 301 -32
rect 244 -46 248 -35
rect 275 -36 301 -33
rect 325 -32 329 -24
rect 313 -36 329 -32
rect 275 -37 306 -36
rect 266 -46 271 -45
rect 275 -46 279 -37
rect 283 -46 287 -45
rect 302 -46 307 -45
rect 325 -46 329 -36
rect 336 -38 340 -34
rect 234 -68 238 -51
rect 293 -68 297 -51
rect 333 -68 337 -51
rect 203 -72 345 -68
rect 119 -89 146 -81
rect -57 -172 -11 -166
rect 123 -246 128 -135
rect 136 -163 146 -89
rect 186 -85 193 -72
rect 283 -76 287 -72
rect 186 -90 280 -85
rect 186 -104 190 -90
rect 211 -104 215 -90
rect 275 -107 280 -90
rect 268 -110 327 -107
rect 167 -131 177 -127
rect 197 -130 201 -113
rect 274 -116 278 -110
rect 282 -130 286 -120
rect 167 -163 171 -131
rect 197 -134 266 -130
rect 282 -133 308 -130
rect 201 -153 205 -149
rect 136 -164 171 -163
rect 136 -168 192 -164
rect 215 -180 220 -134
rect 282 -139 286 -133
rect 186 -215 191 -188
rect 274 -220 278 -143
rect 304 -185 308 -133
rect 324 -169 327 -110
rect 358 -174 365 -7
rect 304 -189 327 -185
rect 191 -225 272 -222
rect 186 -227 272 -225
rect 305 -196 318 -192
rect 305 -246 311 -196
rect 315 -201 318 -196
rect 324 -194 327 -189
rect 324 -198 333 -194
rect 315 -205 347 -201
rect 414 -205 429 -201
rect 123 -251 311 -246
<< m2contact >>
rect 149 22 157 29
rect 10 6 16 12
rect 51 -70 58 -63
rect 119 -35 128 -27
rect -36 -77 -29 -70
rect 141 -72 150 -63
rect 301 -36 306 -31
rect 266 -45 271 -40
rect 283 -45 288 -40
rect 302 -45 307 -40
rect 340 -39 345 -34
rect 91 -95 99 -87
rect 11 -158 19 -151
rect 92 -225 100 -215
rect 51 -232 58 -225
rect 193 -153 201 -146
rect 183 -225 191 -215
rect 272 -227 278 -220
rect 324 -232 330 -226
<< metal2 >>
rect 149 -27 157 22
rect 128 -35 157 -27
rect 317 -30 380 -26
rect 317 -31 322 -30
rect 306 -36 321 -31
rect -69 -47 231 -42
rect 271 -44 283 -40
rect 288 -44 302 -40
rect -36 -70 -29 -66
rect -36 -151 -29 -77
rect -36 -158 11 -151
rect 51 -225 58 -70
rect 91 -72 141 -66
rect 91 -87 98 -72
rect 154 -146 161 -47
rect 227 -61 231 -47
rect 341 -61 345 -39
rect 227 -65 345 -61
rect 154 -153 193 -146
rect 100 -225 183 -216
rect 278 -226 321 -220
rect 278 -227 324 -226
rect 317 -232 324 -227
use 2_input_OR  2_input_OR_0
timestamp 1701467916
transform 1 0 347 0 1 -208
box -23 -24 68 39
use AND  AND_0
timestamp 1700315882
transform 1 0 45 0 1 -136
box -60 -96 78 46
use XOR  XOR_0
timestamp 1701339318
transform 1 0 34 0 1 13
box -20 -32 116 37
<< end >>
