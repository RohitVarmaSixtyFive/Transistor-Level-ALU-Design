magic
tech scmos
timestamp 1701341351
<< nwell >>
rect -23 15 20 32
rect 30 15 65 32
<< ntransistor >>
rect -9 -12 -7 -8
rect 3 -12 5 -8
rect 46 -15 48 -10
<< ptransistor >>
rect -9 22 -7 26
rect 3 22 5 26
rect 46 21 48 26
<< ndiffusion >>
rect -12 -12 -9 -8
rect -7 -12 -4 -8
rect 0 -12 3 -8
rect 5 -12 10 -8
rect 43 -15 46 -10
rect 48 -15 51 -10
<< pdiffusion >>
rect -12 22 -9 26
rect -7 22 3 26
rect 5 22 10 26
rect 43 21 46 26
rect 48 21 51 26
<< ndcontact >>
rect -16 -12 -12 -8
rect -4 -12 0 -8
rect 10 -12 14 -8
rect 38 -15 43 -10
rect 51 -15 56 -10
<< pdcontact >>
rect -16 22 -12 26
rect 10 22 14 26
rect 38 21 43 26
rect 51 21 56 26
<< polysilicon >>
rect -9 26 -7 29
rect 3 26 5 29
rect 46 26 48 29
rect -9 14 -7 22
rect -9 -8 -7 10
rect 3 7 5 22
rect 3 -8 5 3
rect 46 -1 48 21
rect 46 -10 48 -5
rect -9 -16 -7 -12
rect 3 -16 5 -12
rect 46 -18 48 -15
<< polycontact >>
rect -11 10 -7 14
rect 1 3 5 7
rect 44 -5 48 -1
<< metal1 >>
rect -23 33 65 39
rect -16 26 -12 33
rect 38 26 43 33
rect -14 10 -11 14
rect -1 3 1 7
rect 10 -1 14 22
rect 51 7 56 21
rect 51 3 68 7
rect -4 -5 44 -1
rect -4 -8 0 -5
rect 51 -10 56 3
rect -16 -18 -12 -12
rect 10 -18 14 -12
rect 38 -18 43 -15
rect -21 -24 68 -18
<< end >>
