magic
tech scmos
timestamp 1701532374
<< nwell >>
rect 10 -38 64 -11
rect 99 -41 124 -25
rect 9 -189 63 -162
rect 98 -192 123 -176
rect 9 -340 63 -313
rect 98 -343 123 -327
<< ntransistor >>
rect 23 -112 26 -95
rect 36 -112 39 -95
rect 22 -263 25 -246
rect 35 -263 38 -246
rect 22 -414 25 -397
rect 35 -414 38 -397
rect 110 -58 112 -54
rect 109 -209 111 -205
rect 109 -360 111 -356
<< ptransistor >>
rect 22 -31 25 -19
rect 36 -31 39 -19
rect 21 -182 24 -170
rect 35 -182 38 -170
rect 21 -333 24 -321
rect 35 -333 38 -321
rect 110 -35 112 -31
rect 109 -186 111 -182
rect 109 -337 111 -333
<< ndiffusion >>
rect 15 -103 17 -95
rect 22 -103 23 -95
rect 15 -112 23 -103
rect 26 -112 36 -95
rect 39 -103 46 -95
rect 51 -103 53 -95
rect 39 -112 53 -103
rect 14 -254 16 -246
rect 21 -254 22 -246
rect 14 -263 22 -254
rect 25 -263 35 -246
rect 38 -254 45 -246
rect 50 -254 52 -246
rect 38 -263 52 -254
rect 14 -405 16 -397
rect 21 -405 22 -397
rect 14 -414 22 -405
rect 25 -414 35 -397
rect 38 -405 45 -397
rect 50 -405 52 -397
rect 38 -414 52 -405
rect 109 -58 110 -54
rect 112 -58 113 -54
rect 108 -209 109 -205
rect 111 -209 112 -205
rect 108 -360 109 -356
rect 111 -360 112 -356
<< pdiffusion >>
rect 16 -28 17 -19
rect 21 -28 22 -19
rect 16 -31 22 -28
rect 25 -28 28 -19
rect 32 -28 36 -19
rect 25 -31 36 -28
rect 39 -28 42 -19
rect 46 -28 49 -19
rect 39 -31 49 -28
rect 15 -179 16 -170
rect 20 -179 21 -170
rect 15 -182 21 -179
rect 24 -179 27 -170
rect 31 -179 35 -170
rect 24 -182 35 -179
rect 38 -179 41 -170
rect 45 -179 48 -170
rect 38 -182 48 -179
rect 15 -330 16 -321
rect 20 -330 21 -321
rect 15 -333 21 -330
rect 24 -330 27 -321
rect 31 -330 35 -321
rect 24 -333 35 -330
rect 38 -330 41 -321
rect 45 -330 48 -321
rect 38 -333 48 -330
rect 109 -35 110 -31
rect 112 -35 113 -31
rect 108 -186 109 -182
rect 111 -186 112 -182
rect 108 -337 109 -333
rect 111 -337 112 -333
<< ndcontact >>
rect 17 -103 22 -95
rect 46 -103 51 -95
rect 16 -254 21 -246
rect 45 -254 50 -246
rect 16 -405 21 -397
rect 45 -405 50 -397
rect 105 -58 109 -54
rect 113 -58 117 -54
rect 104 -209 108 -205
rect 112 -209 116 -205
rect 104 -360 108 -356
rect 112 -360 116 -356
<< pdcontact >>
rect 17 -28 21 -19
rect 28 -28 32 -19
rect 42 -28 46 -19
rect 16 -179 20 -170
rect 27 -179 31 -170
rect 41 -179 45 -170
rect 16 -330 20 -321
rect 27 -330 31 -321
rect 41 -330 45 -321
rect 105 -35 109 -31
rect 113 -35 117 -31
rect 104 -186 108 -182
rect 112 -186 116 -182
rect 104 -337 108 -333
rect 112 -337 116 -333
<< polysilicon >>
rect 74 1 78 143
rect 22 -19 25 -9
rect 36 -19 39 -8
rect 22 -43 25 -31
rect 12 -46 25 -43
rect 36 -64 39 -31
rect 23 -95 26 -83
rect 36 -95 39 -68
rect 23 -116 26 -112
rect 36 -116 39 -112
rect 74 -150 78 -5
rect 21 -170 24 -160
rect 35 -170 38 -159
rect 21 -194 24 -182
rect 11 -197 24 -194
rect 35 -215 38 -182
rect 22 -246 25 -234
rect 35 -246 38 -219
rect 22 -267 25 -263
rect 35 -267 38 -263
rect 74 -301 78 -156
rect 21 -321 24 -311
rect 35 -321 38 -310
rect 21 -345 24 -333
rect 11 -348 24 -345
rect 35 -366 38 -333
rect 22 -397 25 -385
rect 35 -397 38 -370
rect 22 -418 25 -414
rect 35 -418 38 -414
rect 74 -445 78 -307
rect 85 -136 89 6
rect 110 -31 112 -28
rect 110 -46 112 -35
rect 101 -49 112 -46
rect 110 -54 112 -49
rect 110 -61 112 -58
rect 85 -287 89 -142
rect 109 -182 111 -179
rect 109 -197 111 -186
rect 100 -200 111 -197
rect 109 -205 111 -200
rect 109 -212 111 -209
rect 85 -438 89 -293
rect 109 -333 111 -330
rect 109 -348 111 -337
rect 100 -351 111 -348
rect 109 -356 111 -351
rect 109 -363 111 -360
rect 85 -445 89 -444
<< polycontact >>
rect 72 143 78 149
rect 72 -5 78 1
rect 8 -46 12 -42
rect 36 -68 40 -64
rect 23 -83 27 -79
rect 72 -156 78 -150
rect 7 -197 11 -193
rect 35 -219 39 -215
rect 22 -234 26 -230
rect 72 -307 78 -301
rect 7 -348 11 -344
rect 35 -370 39 -366
rect 22 -385 26 -381
rect 85 6 91 12
rect 97 -49 101 -45
rect 85 -142 91 -136
rect 96 -200 100 -196
rect 85 -293 91 -287
rect 96 -351 100 -347
rect 85 -444 91 -438
<< metal1 >>
rect 56 146 64 157
rect 135 100 147 103
rect -7 95 2 99
rect 21 80 32 84
rect 56 4 61 9
rect 17 -5 72 0
rect 78 -5 111 0
rect 17 -19 21 -5
rect 42 -19 46 -5
rect 106 -22 111 -5
rect 99 -25 124 -22
rect -2 -46 8 -42
rect 28 -45 32 -28
rect 105 -31 109 -25
rect 113 -45 117 -35
rect -2 -79 2 -46
rect 28 -49 97 -45
rect 113 -48 147 -45
rect 29 -68 36 -64
rect -2 -83 23 -79
rect 46 -95 51 -49
rect 113 -54 117 -48
rect 17 -137 22 -103
rect 17 -142 85 -137
rect 105 -137 109 -58
rect 91 -142 109 -137
rect 16 -156 72 -151
rect 78 -156 110 -151
rect 16 -170 20 -156
rect 41 -170 45 -156
rect 105 -173 110 -156
rect 98 -176 123 -173
rect -3 -197 7 -193
rect 27 -196 31 -179
rect 104 -182 108 -176
rect 112 -196 116 -186
rect -3 -230 1 -197
rect 27 -200 96 -196
rect 112 -199 144 -196
rect 28 -219 35 -215
rect -3 -234 22 -230
rect 45 -246 50 -200
rect 112 -205 116 -199
rect 16 -288 21 -254
rect 16 -293 85 -288
rect 104 -288 108 -209
rect 91 -293 108 -288
rect 16 -307 72 -302
rect 78 -307 110 -302
rect 16 -321 20 -307
rect 41 -321 45 -307
rect 105 -324 110 -307
rect 98 -327 123 -324
rect -3 -348 7 -344
rect 27 -347 31 -330
rect 104 -333 108 -327
rect 112 -347 116 -337
rect -3 -381 1 -348
rect 27 -351 96 -347
rect 112 -350 145 -347
rect 28 -370 35 -366
rect -3 -385 22 -381
rect 45 -397 50 -351
rect 112 -356 116 -350
rect 16 -439 21 -405
rect 16 -444 85 -439
rect 104 -439 108 -360
rect 91 -444 108 -439
use AND  AND_0
timestamp 1700315882
transform 1 0 58 0 1 102
box -60 -96 78 46
<< labels >>
rlabel metal1 -1 -54 1 -52 3 a1
rlabel metal1 -2 -207 0 -205 3 a2
rlabel metal1 -2 -356 0 -354 3 a3
rlabel metal1 29 -369 31 -367 1 b3
rlabel metal1 30 -218 32 -216 1 b2
rlabel metal1 30 -67 32 -65 1 b1
rlabel metal1 145 101 146 102 7 and_out0
rlabel metal1 143 -47 144 -46 7 and_out1
rlabel metal1 140 -198 141 -197 1 and_out2
rlabel metal1 142 -349 143 -348 7 and_out3
rlabel metal1 -7 96 -5 98 3 a0
rlabel metal1 22 81 24 82 1 b0
<< end >>
