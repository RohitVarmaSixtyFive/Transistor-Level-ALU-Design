magic
tech scmos
timestamp 1699298635
<< nwell >>
rect 66 21 124 22
rect -30 3 30 20
rect 66 4 125 21
<< ntransistor >>
rect -18 -31 -16 -27
rect -7 -31 -5 -27
rect 5 -31 7 -27
rect 15 -31 17 -27
rect 94 -34 96 -28
<< ptransistor >>
rect -18 9 -16 13
rect -7 9 -5 13
rect 5 9 7 13
rect 15 9 17 13
rect 94 10 96 16
<< ndiffusion >>
rect -19 -31 -18 -27
rect -16 -31 -13 -27
rect -9 -31 -7 -27
rect -5 -31 -2 -27
rect 2 -31 5 -27
rect 7 -31 9 -27
rect 13 -31 15 -27
rect 17 -31 20 -27
rect 90 -34 94 -28
rect 96 -34 99 -28
<< pdiffusion >>
rect -19 9 -18 13
rect -16 9 -7 13
rect -5 9 5 13
rect 7 9 15 13
rect 17 9 18 13
rect 91 10 94 16
rect 96 10 99 16
<< ndcontact >>
rect -23 -31 -19 -27
rect -13 -31 -9 -27
rect -2 -31 2 -27
rect 9 -31 13 -27
rect 20 -31 24 -27
rect 86 -34 90 -28
rect 99 -34 103 -28
<< pdcontact >>
rect -23 9 -19 13
rect 18 9 22 13
rect 86 10 91 16
rect 99 10 103 16
<< polysilicon >>
rect -18 13 -16 16
rect -7 13 -5 17
rect 5 13 7 17
rect 15 13 17 17
rect 94 16 96 20
rect -18 2 -16 9
rect -29 -2 -16 2
rect -7 -4 -5 9
rect 5 -1 7 9
rect 15 2 17 9
rect 15 -1 20 2
rect 94 -3 96 10
rect -30 -15 -16 -11
rect -18 -27 -16 -15
rect -7 -27 -5 -8
rect 5 -27 7 -5
rect 15 -15 20 -12
rect 15 -27 17 -15
rect 94 -28 96 -8
rect -18 -39 -16 -31
rect -7 -38 -5 -31
rect 5 -39 7 -31
rect 15 -38 17 -31
rect 94 -40 96 -34
<< polycontact >>
rect -35 -2 -29 2
rect -9 -8 -5 -4
rect 3 -5 7 -1
rect 20 -2 24 2
rect -36 -15 -30 -11
rect 84 -8 96 -3
rect 20 -15 24 -11
<< metal1 >>
rect -30 22 127 28
rect -30 20 38 22
rect -23 13 -19 20
rect 86 16 91 22
rect 22 9 33 13
rect -44 -2 -35 2
rect -44 -11 -41 -2
rect -12 -8 -9 -4
rect 0 -5 3 -1
rect 20 -11 24 -2
rect -44 -15 -36 -11
rect 29 -3 33 9
rect 29 -8 84 -3
rect 99 -8 103 10
rect 29 -20 33 -8
rect -23 -23 33 -20
rect 99 -14 114 -8
rect -23 -27 -19 -23
rect -2 -27 2 -23
rect 20 -27 24 -23
rect 99 -28 103 -14
rect -13 -37 -9 -31
rect 9 -37 13 -31
rect 86 -37 90 -34
rect -25 -46 114 -37
rect -25 -48 85 -46
<< labels >>
rlabel metal1 9 23 12 24 5 VDD
rlabel metal1 -38 -1 -37 0 1 a
rlabel metal1 -10 -7 -9 -6 1 b
rlabel metal1 2 -4 3 -3 1 c
rlabel metal1 22 -7 23 -6 1 d
rlabel metal1 52 -45 55 -43 1 gnd
rlabel metal1 79 -6 80 -5 1 in
rlabel metal1 108 -12 109 -11 1 out
<< end >>
