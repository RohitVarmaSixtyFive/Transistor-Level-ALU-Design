magic
tech scmos
timestamp 1701545594
<< nwell >>
rect 213 -406 324 -379
rect 391 -392 416 -376
rect 232 -584 335 -557
rect 374 -570 399 -554
rect 525 -664 585 -647
rect 621 -665 680 -648
rect 621 -666 679 -665
rect 252 -747 334 -720
rect 341 -733 366 -717
rect 251 -915 305 -888
rect 340 -901 365 -885
<< ntransistor >>
rect 226 -322 229 -305
rect 247 -322 250 -305
rect 269 -322 272 -305
rect 293 -322 296 -305
rect 315 -322 318 -305
rect 402 -363 404 -359
rect 245 -500 248 -483
rect 266 -500 269 -483
rect 288 -500 291 -483
rect 312 -500 315 -483
rect 385 -541 387 -537
rect 265 -663 268 -646
rect 286 -663 289 -646
rect 308 -663 311 -646
rect 537 -617 539 -613
rect 548 -617 550 -613
rect 560 -617 562 -613
rect 570 -617 572 -613
rect 649 -616 651 -610
rect 352 -704 354 -700
rect 264 -831 267 -814
rect 277 -831 280 -814
rect 351 -872 353 -868
<< ptransistor >>
rect 225 -398 228 -386
rect 247 -398 250 -386
rect 267 -398 270 -386
rect 287 -398 290 -386
rect 307 -398 310 -386
rect 402 -386 404 -382
rect 244 -576 247 -564
rect 266 -576 269 -564
rect 286 -576 289 -564
rect 306 -576 309 -564
rect 385 -564 387 -560
rect 537 -657 539 -653
rect 548 -657 550 -653
rect 560 -657 562 -653
rect 570 -657 572 -653
rect 649 -660 651 -654
rect 264 -739 267 -727
rect 286 -739 289 -727
rect 306 -739 309 -727
rect 352 -727 354 -723
rect 351 -895 353 -891
rect 263 -907 266 -895
rect 277 -907 280 -895
<< ndiffusion >>
rect 218 -314 226 -305
rect 218 -322 220 -314
rect 225 -322 226 -314
rect 229 -322 247 -305
rect 250 -322 269 -305
rect 272 -322 293 -305
rect 296 -322 315 -305
rect 318 -314 326 -305
rect 318 -322 320 -314
rect 325 -322 326 -314
rect 401 -363 402 -359
rect 404 -363 405 -359
rect 237 -492 245 -483
rect 237 -500 239 -492
rect 244 -500 245 -492
rect 248 -500 266 -483
rect 269 -500 288 -483
rect 291 -500 312 -483
rect 315 -493 325 -483
rect 315 -500 320 -493
rect 384 -541 385 -537
rect 387 -541 388 -537
rect 257 -655 265 -646
rect 257 -663 259 -655
rect 264 -663 265 -655
rect 268 -663 286 -646
rect 289 -663 308 -646
rect 311 -654 326 -646
rect 311 -663 320 -654
rect 536 -617 537 -613
rect 539 -617 542 -613
rect 546 -617 548 -613
rect 550 -617 553 -613
rect 557 -617 560 -613
rect 562 -617 564 -613
rect 568 -617 570 -613
rect 572 -617 575 -613
rect 645 -616 649 -610
rect 651 -616 654 -610
rect 351 -704 352 -700
rect 354 -704 355 -700
rect 256 -823 264 -814
rect 256 -831 258 -823
rect 263 -831 264 -823
rect 267 -831 277 -814
rect 280 -823 294 -814
rect 280 -831 287 -823
rect 292 -831 294 -823
rect 350 -872 351 -868
rect 353 -872 354 -868
<< pdiffusion >>
rect 219 -389 225 -386
rect 219 -398 220 -389
rect 224 -398 225 -389
rect 228 -389 247 -386
rect 228 -398 234 -389
rect 238 -398 247 -389
rect 250 -389 267 -386
rect 250 -398 256 -389
rect 260 -398 267 -389
rect 270 -389 287 -386
rect 270 -398 275 -389
rect 279 -398 287 -389
rect 290 -389 307 -386
rect 290 -398 299 -389
rect 303 -398 307 -389
rect 310 -389 318 -386
rect 310 -398 311 -389
rect 315 -398 318 -389
rect 401 -386 402 -382
rect 404 -386 405 -382
rect 238 -567 244 -564
rect 238 -576 239 -567
rect 243 -576 244 -567
rect 247 -567 266 -564
rect 247 -576 253 -567
rect 257 -576 266 -567
rect 269 -567 286 -564
rect 269 -576 275 -567
rect 279 -576 286 -567
rect 289 -567 306 -564
rect 289 -576 294 -567
rect 298 -576 306 -567
rect 309 -567 325 -564
rect 309 -576 318 -567
rect 322 -576 325 -567
rect 384 -564 385 -560
rect 387 -564 388 -560
rect 536 -657 537 -653
rect 539 -657 548 -653
rect 550 -657 560 -653
rect 562 -657 570 -653
rect 572 -657 573 -653
rect 646 -660 649 -654
rect 651 -660 654 -654
rect 258 -730 264 -727
rect 258 -739 259 -730
rect 263 -739 264 -730
rect 267 -730 286 -727
rect 267 -739 273 -730
rect 277 -739 286 -730
rect 289 -730 306 -727
rect 289 -739 295 -730
rect 299 -739 306 -730
rect 309 -730 326 -727
rect 309 -739 314 -730
rect 318 -739 326 -730
rect 351 -727 352 -723
rect 354 -727 355 -723
rect 350 -895 351 -891
rect 353 -895 354 -891
rect 257 -898 263 -895
rect 257 -907 258 -898
rect 262 -907 263 -898
rect 266 -898 277 -895
rect 266 -907 269 -898
rect 273 -907 277 -898
rect 280 -898 290 -895
rect 280 -907 283 -898
rect 287 -907 290 -898
<< ndcontact >>
rect 220 -322 225 -314
rect 320 -322 325 -314
rect 397 -363 401 -359
rect 405 -363 409 -359
rect 239 -500 244 -492
rect 320 -500 325 -493
rect 380 -541 384 -537
rect 388 -541 392 -537
rect 259 -663 264 -655
rect 320 -663 326 -654
rect 532 -617 536 -613
rect 542 -617 546 -613
rect 553 -617 557 -613
rect 564 -617 568 -613
rect 575 -617 579 -613
rect 641 -616 645 -610
rect 654 -616 658 -610
rect 347 -704 351 -700
rect 355 -704 359 -700
rect 258 -831 263 -823
rect 287 -831 292 -823
rect 346 -872 350 -868
rect 354 -872 358 -868
<< pdcontact >>
rect 220 -398 224 -389
rect 234 -398 238 -389
rect 256 -398 260 -389
rect 275 -398 279 -389
rect 299 -398 303 -389
rect 311 -398 315 -389
rect 397 -386 401 -382
rect 405 -386 409 -382
rect 239 -576 243 -567
rect 253 -576 257 -567
rect 275 -576 279 -567
rect 294 -576 298 -567
rect 318 -576 322 -567
rect 380 -564 384 -560
rect 388 -564 392 -560
rect 532 -657 536 -653
rect 573 -657 577 -653
rect 641 -660 646 -654
rect 654 -660 658 -654
rect 259 -739 263 -730
rect 273 -739 277 -730
rect 295 -739 299 -730
rect 314 -739 318 -730
rect 347 -727 351 -723
rect 355 -727 359 -723
rect 346 -895 350 -891
rect 354 -895 358 -891
rect 258 -907 262 -898
rect 269 -907 273 -898
rect 283 -907 287 -898
<< polysilicon >>
rect 355 752 398 760
rect 333 566 340 626
rect 390 600 398 752
rect 390 597 599 600
rect 356 592 599 597
rect 356 589 398 592
rect 324 559 340 566
rect 324 521 331 559
rect 390 534 398 589
rect 378 526 398 534
rect 324 514 339 521
rect 332 465 339 514
rect 332 456 339 459
rect 332 451 360 456
rect 354 304 360 451
rect 378 437 386 526
rect 591 517 599 592
rect 386 428 435 436
rect 427 361 435 428
rect 537 423 544 436
rect 396 353 435 361
rect 501 416 544 423
rect 82 204 235 206
rect -54 88 31 90
rect -54 -362 -52 88
rect -2 81 3 82
rect -21 1 -17 2
rect -47 -3 -17 1
rect -47 -350 -43 -3
rect -2 -8 3 77
rect 27 73 31 88
rect 82 72 84 204
rect 354 123 360 295
rect 396 265 404 353
rect 395 264 467 265
rect 404 254 467 264
rect 412 114 430 124
rect 117 82 122 83
rect 117 77 327 82
rect 14 -3 31 2
rect -2 -98 3 -12
rect 27 -16 31 -3
rect 82 -17 84 -5
rect 112 -73 116 12
rect 322 -17 327 77
rect 116 -77 208 -73
rect -14 -350 -11 -183
rect -2 -187 3 -102
rect 26 -84 30 -83
rect 26 -86 102 -84
rect 26 -106 30 -86
rect 81 -106 83 -94
rect 112 -163 116 -77
rect 128 -85 137 -83
rect 135 -96 137 -85
rect 26 -194 30 -183
rect 81 -195 83 -183
rect 112 -252 116 -167
rect 129 -98 137 -96
rect 129 -362 131 -98
rect 204 -155 208 -77
rect 424 -154 430 114
rect 459 -9 467 254
rect 459 -14 468 -9
rect 204 -159 319 -155
rect 424 -272 430 -160
rect 440 -16 468 -14
rect 440 -22 460 -16
rect 440 -165 448 -22
rect 501 -92 508 416
rect 470 -99 508 -92
rect 440 -173 467 -165
rect 226 -305 229 -301
rect 247 -305 250 -301
rect 269 -305 272 -301
rect 293 -305 296 -301
rect 315 -305 318 -301
rect 226 -334 229 -322
rect 247 -342 250 -322
rect 269 -342 272 -322
rect 293 -342 296 -322
rect 315 -343 318 -322
rect 317 -347 318 -343
rect -54 -364 235 -362
rect -14 -385 -10 -383
rect -12 -850 -10 -385
rect 129 -427 131 -364
rect 215 -374 228 -371
rect 225 -386 228 -374
rect 247 -386 250 -363
rect 267 -386 270 -363
rect 287 -386 290 -363
rect 313 -374 317 -363
rect 307 -377 317 -374
rect 307 -386 310 -377
rect 225 -408 228 -398
rect 247 -409 250 -398
rect 267 -408 270 -398
rect 287 -409 290 -398
rect 307 -409 310 -398
rect 113 -429 131 -427
rect 113 -683 115 -429
rect 354 -453 360 -281
rect 412 -282 430 -272
rect 402 -359 404 -356
rect 402 -368 404 -363
rect 393 -371 404 -368
rect 402 -382 404 -371
rect 402 -389 404 -386
rect 459 -412 467 -173
rect 404 -422 467 -412
rect 395 -423 467 -422
rect 245 -483 248 -479
rect 266 -483 269 -479
rect 288 -483 291 -479
rect 312 -483 315 -479
rect 245 -512 248 -500
rect 266 -520 269 -500
rect 288 -520 291 -500
rect 312 -520 315 -500
rect 234 -552 247 -549
rect 244 -564 247 -552
rect 266 -564 269 -541
rect 286 -564 289 -541
rect 306 -564 309 -541
rect 244 -586 247 -576
rect 266 -587 269 -576
rect 286 -586 289 -576
rect 306 -587 309 -576
rect 354 -609 360 -462
rect 396 -511 404 -423
rect 396 -519 435 -511
rect 385 -537 387 -534
rect 385 -546 387 -541
rect 376 -549 387 -546
rect 385 -560 387 -549
rect 385 -567 387 -564
rect 427 -586 435 -519
rect 501 -574 508 -99
rect 501 -581 544 -574
rect 332 -614 360 -609
rect 386 -594 435 -586
rect 537 -594 544 -581
rect 332 -617 339 -614
rect 265 -646 268 -642
rect 286 -646 289 -642
rect 308 -646 311 -642
rect 265 -675 268 -663
rect 286 -683 289 -663
rect 308 -683 311 -663
rect 332 -672 339 -623
rect 324 -679 339 -672
rect 113 -686 286 -683
rect 274 -687 286 -686
rect 254 -715 267 -712
rect 264 -727 267 -715
rect 286 -727 289 -704
rect 306 -727 309 -704
rect 324 -717 331 -679
rect 378 -684 386 -595
rect 537 -613 539 -605
rect 548 -613 550 -606
rect 560 -613 562 -605
rect 570 -613 572 -606
rect 649 -610 651 -604
rect 537 -629 539 -617
rect 525 -633 539 -629
rect 548 -636 550 -617
rect 560 -639 562 -617
rect 570 -629 572 -617
rect 570 -632 575 -629
rect 649 -636 651 -616
rect 526 -646 539 -642
rect 537 -653 539 -646
rect 548 -653 550 -640
rect 560 -653 562 -643
rect 570 -646 575 -643
rect 570 -653 572 -646
rect 649 -654 651 -641
rect 537 -660 539 -657
rect 548 -661 550 -657
rect 560 -661 562 -657
rect 570 -661 572 -657
rect 649 -664 651 -660
rect 378 -692 398 -684
rect 352 -700 354 -697
rect 352 -709 354 -704
rect 343 -712 354 -709
rect 324 -724 340 -717
rect 352 -723 354 -712
rect 264 -749 267 -739
rect 286 -750 289 -739
rect 306 -749 309 -739
rect 333 -784 340 -724
rect 352 -730 354 -727
rect 390 -747 398 -692
rect 356 -750 398 -747
rect 591 -750 599 -675
rect 356 -755 599 -750
rect 390 -758 599 -755
rect 264 -814 267 -810
rect 277 -814 280 -810
rect 264 -843 267 -831
rect -12 -852 196 -850
rect 277 -858 280 -831
rect 253 -883 266 -880
rect 263 -895 266 -883
rect 277 -895 280 -862
rect 351 -868 353 -865
rect 351 -877 353 -872
rect 342 -880 353 -877
rect 351 -891 353 -880
rect 351 -898 353 -895
rect 263 -917 266 -907
rect 277 -918 280 -907
rect 390 -910 398 -758
rect 355 -918 398 -910
<< polycontact >>
rect 347 752 355 760
rect 333 626 340 632
rect 348 589 356 597
rect 332 459 339 465
rect 591 507 601 517
rect 378 428 386 437
rect 537 436 544 442
rect 354 295 363 304
rect -2 77 3 81
rect -17 -3 -12 2
rect 235 203 239 207
rect 395 254 404 264
rect 354 114 363 123
rect 400 114 412 124
rect 111 77 117 83
rect 112 12 116 16
rect 9 -3 14 2
rect -2 -12 3 -8
rect 82 -5 86 -1
rect 322 -24 329 -17
rect 112 -77 116 -73
rect -2 -102 3 -98
rect -15 -183 -9 -177
rect 102 -86 106 -82
rect 81 -94 85 -90
rect 124 -86 128 -82
rect 112 -167 116 -163
rect 24 -183 30 -177
rect -2 -191 3 -187
rect 81 -183 86 -178
rect 112 -256 116 -252
rect -47 -356 -41 -350
rect -15 -355 -9 -350
rect 319 -160 326 -154
rect 424 -160 430 -154
rect 460 -24 468 -16
rect 461 -99 470 -91
rect 354 -281 363 -272
rect 226 -338 230 -334
rect 247 -346 251 -342
rect 269 -346 273 -342
rect 292 -346 296 -342
rect 313 -347 317 -343
rect -15 -383 -9 -378
rect 235 -365 239 -361
rect 247 -363 251 -359
rect 266 -363 270 -359
rect 211 -375 215 -371
rect 287 -363 291 -359
rect 313 -363 317 -359
rect 400 -282 412 -272
rect 389 -372 393 -368
rect 395 -422 404 -412
rect 354 -462 363 -453
rect 245 -516 249 -512
rect 266 -524 270 -520
rect 288 -524 292 -520
rect 311 -524 315 -520
rect 266 -541 270 -537
rect 285 -541 289 -537
rect 230 -553 234 -549
rect 306 -541 310 -537
rect 372 -550 376 -546
rect 378 -595 386 -586
rect 332 -623 339 -617
rect 265 -679 269 -675
rect 286 -687 290 -683
rect 308 -687 312 -683
rect 286 -704 290 -700
rect 305 -704 309 -700
rect 250 -716 254 -712
rect 537 -600 544 -594
rect 519 -633 525 -629
rect 546 -640 550 -636
rect 575 -633 579 -629
rect 520 -646 526 -642
rect 558 -643 562 -639
rect 639 -641 651 -636
rect 575 -646 579 -642
rect 591 -675 601 -665
rect 339 -713 343 -709
rect 348 -755 356 -747
rect 333 -790 340 -784
rect 264 -847 268 -843
rect 196 -853 202 -848
rect 277 -862 281 -858
rect 249 -884 253 -880
rect 338 -881 342 -877
rect 347 -918 355 -910
<< metal1 >>
rect -61 715 -57 717
rect -61 711 211 715
rect -61 -216 -57 711
rect 151 690 243 695
rect -43 542 105 546
rect -43 -127 -39 542
rect -28 394 103 398
rect -28 -37 -24 394
rect -17 213 110 217
rect -17 52 -13 213
rect 51 80 55 86
rect -17 48 -4 52
rect 51 7 56 13
rect -12 -3 9 2
rect 14 -3 15 2
rect 120 -1 124 375
rect 86 -5 125 -1
rect -28 -41 -4 -37
rect 106 -86 124 -82
rect 139 -90 143 526
rect 85 -94 143 -90
rect -43 -131 -5 -127
rect -9 -183 24 -177
rect 151 -178 156 690
rect 493 544 498 565
rect 184 521 189 524
rect 163 -24 168 194
rect 174 192 177 367
rect 162 -29 168 -24
rect 172 190 177 192
rect 172 -120 177 185
rect 184 363 189 515
rect 553 481 556 485
rect 571 478 579 481
rect 184 181 189 357
rect 510 214 513 475
rect 666 472 713 478
rect 422 211 513 214
rect 86 -183 156 -178
rect 184 -199 189 174
rect 483 -67 609 -64
rect 224 -83 230 -80
rect 133 -204 189 -199
rect 194 -129 200 -125
rect 133 -208 139 -204
rect -62 -220 -5 -216
rect 194 -220 198 -129
rect 161 -225 198 -220
rect -47 -554 -41 -356
rect -28 -383 -22 -359
rect -15 -378 -9 -355
rect -2 -395 4 -357
rect 132 -382 138 -349
rect 161 -352 166 -225
rect 226 -235 229 -83
rect 186 -238 229 -235
rect 186 -332 189 -238
rect 220 -280 354 -272
rect 220 -314 225 -280
rect 363 -280 400 -272
rect 398 -282 400 -280
rect 201 -338 226 -334
rect 161 -357 193 -352
rect -36 -401 4 -395
rect -36 -534 -30 -401
rect 161 -514 166 -357
rect 201 -371 205 -338
rect 235 -346 247 -342
rect 256 -346 269 -342
rect 280 -343 292 -342
rect 235 -359 240 -346
rect 256 -352 261 -346
rect 256 -359 261 -357
rect 286 -346 292 -343
rect 280 -359 285 -348
rect 308 -347 313 -343
rect 300 -359 305 -350
rect 235 -361 247 -359
rect 239 -363 247 -361
rect 256 -363 266 -359
rect 280 -363 287 -359
rect 300 -363 313 -359
rect 320 -369 325 -322
rect 398 -350 404 -282
rect 391 -355 410 -350
rect 397 -359 401 -355
rect 206 -375 211 -371
rect 234 -372 389 -369
rect 234 -373 393 -372
rect 405 -369 409 -363
rect 405 -372 513 -369
rect 234 -389 238 -373
rect 275 -389 279 -373
rect 311 -389 315 -373
rect 405 -382 409 -372
rect 397 -392 401 -386
rect 391 -395 416 -392
rect 220 -412 224 -398
rect 256 -412 260 -398
rect 299 -412 303 -398
rect 398 -412 403 -395
rect 220 -417 395 -412
rect 239 -458 354 -454
rect 239 -492 244 -458
rect 363 -458 387 -454
rect 161 -519 196 -514
rect 220 -516 245 -512
rect -36 -541 -26 -534
rect 129 -547 137 -532
rect 220 -549 224 -516
rect 254 -524 266 -520
rect 275 -524 288 -520
rect 306 -523 311 -520
rect 299 -524 311 -523
rect 254 -534 259 -524
rect 275 -525 280 -524
rect 275 -537 280 -530
rect 299 -537 304 -524
rect 259 -541 266 -537
rect 275 -541 285 -537
rect 299 -541 306 -537
rect 320 -546 325 -500
rect 381 -528 387 -458
rect 374 -533 393 -528
rect 380 -537 384 -533
rect 217 -553 230 -549
rect 253 -550 372 -546
rect 388 -547 392 -541
rect 388 -550 405 -547
rect 217 -554 223 -553
rect -47 -560 102 -554
rect 96 -569 102 -560
rect 160 -560 223 -554
rect 160 -569 166 -560
rect 253 -567 257 -550
rect 294 -567 298 -550
rect 388 -560 392 -550
rect 96 -575 166 -569
rect 380 -570 384 -564
rect 374 -573 399 -570
rect -25 -668 -17 -585
rect 239 -590 243 -576
rect 275 -590 279 -576
rect 318 -590 322 -576
rect 381 -586 386 -573
rect 239 -595 378 -590
rect 259 -621 332 -617
rect 259 -655 264 -621
rect 339 -621 354 -617
rect -25 -676 194 -668
rect 240 -679 265 -675
rect 240 -700 244 -679
rect 274 -687 286 -683
rect 302 -687 308 -683
rect 274 -700 279 -687
rect 295 -700 300 -687
rect 274 -704 286 -700
rect 295 -704 305 -700
rect 240 -712 244 -707
rect 320 -709 326 -663
rect 348 -691 354 -621
rect 510 -629 513 -372
rect 530 -600 537 -596
rect 544 -598 640 -596
rect 544 -600 669 -598
rect 530 -607 669 -600
rect 542 -613 546 -607
rect 564 -613 568 -607
rect 641 -610 645 -607
rect 532 -621 536 -617
rect 553 -621 557 -617
rect 575 -621 579 -617
rect 532 -624 588 -621
rect 510 -633 519 -629
rect 511 -642 514 -633
rect 575 -636 579 -633
rect 544 -640 546 -636
rect 511 -646 520 -642
rect 553 -643 558 -639
rect 571 -639 579 -636
rect 575 -642 579 -639
rect 584 -636 588 -624
rect 654 -630 658 -616
rect 654 -636 713 -630
rect 584 -641 639 -636
rect 584 -653 588 -641
rect 577 -657 588 -653
rect 654 -654 658 -636
rect 532 -664 536 -657
rect 525 -665 593 -664
rect 525 -672 591 -665
rect 641 -666 646 -660
rect 601 -672 682 -666
rect 341 -696 360 -691
rect 347 -700 351 -696
rect 240 -716 250 -712
rect 273 -713 339 -709
rect 355 -710 359 -704
rect 355 -713 381 -710
rect 273 -730 277 -713
rect 314 -730 318 -713
rect 355 -723 359 -713
rect 493 -723 498 -702
rect 347 -733 351 -727
rect 341 -736 366 -733
rect 259 -753 263 -739
rect 295 -753 299 -739
rect 348 -747 353 -736
rect 259 -755 348 -753
rect 259 -758 353 -755
rect 258 -789 333 -784
rect 258 -823 263 -789
rect 340 -789 350 -784
rect 239 -847 264 -843
rect 239 -848 243 -847
rect 202 -853 243 -848
rect 239 -880 243 -853
rect 271 -862 277 -858
rect 287 -877 292 -831
rect 346 -868 350 -789
rect 239 -884 249 -880
rect 269 -881 338 -877
rect 354 -878 358 -872
rect 354 -881 376 -878
rect 269 -898 273 -881
rect 354 -891 358 -881
rect 346 -901 350 -895
rect 340 -904 365 -901
rect 258 -921 262 -907
rect 283 -921 287 -907
rect 347 -910 352 -904
rect 347 -921 352 -918
rect 258 -926 352 -921
<< m2contact >>
rect 376 720 381 725
rect 211 711 219 719
rect 260 700 271 708
rect 105 542 113 549
rect 134 526 143 534
rect 103 394 109 400
rect 120 375 127 382
rect 110 213 116 219
rect 492 565 499 571
rect 381 552 386 557
rect 237 542 245 549
rect 492 538 499 544
rect 270 526 279 535
rect 295 523 302 529
rect 184 515 191 521
rect 174 367 180 372
rect 163 194 169 199
rect 162 -35 168 -29
rect 172 185 177 190
rect 172 -125 177 -120
rect 552 485 557 490
rect 539 478 544 483
rect 566 478 571 483
rect 218 394 224 400
rect 405 389 410 394
rect 251 376 259 383
rect 275 367 280 372
rect 184 357 191 363
rect 299 358 306 365
rect 201 213 206 218
rect 255 194 261 199
rect 280 185 286 190
rect 300 185 308 192
rect 184 174 191 181
rect 224 -80 230 -74
rect 354 -82 360 -76
rect 194 -125 200 -119
rect 133 -214 139 -208
rect 132 -349 138 -342
rect -28 -359 -22 -353
rect -2 -357 4 -351
rect -28 -389 -22 -383
rect 132 -389 138 -382
rect 378 -84 384 -78
rect 333 -90 339 -84
rect 298 -100 304 -94
rect 186 -339 192 -332
rect 193 -357 198 -352
rect 255 -357 261 -352
rect 280 -348 286 -343
rect 300 -350 308 -343
rect 201 -376 206 -371
rect 196 -520 204 -513
rect -26 -541 -16 -531
rect 129 -532 137 -525
rect 129 -554 137 -547
rect 299 -523 306 -516
rect 251 -541 259 -534
rect 275 -530 280 -525
rect 405 -552 410 -547
rect -26 -585 -16 -575
rect 194 -679 205 -668
rect 295 -687 302 -681
rect 237 -707 245 -700
rect 539 -641 544 -636
rect 566 -641 571 -636
rect 552 -648 557 -643
rect 492 -702 499 -696
rect 381 -715 386 -710
rect 492 -729 499 -723
rect 260 -866 271 -858
rect 376 -883 381 -878
<< metal2 >>
rect 381 720 498 725
rect 219 711 265 719
rect 260 708 265 711
rect 493 571 498 720
rect 388 557 557 558
rect 386 553 557 557
rect 386 552 391 553
rect 113 542 237 549
rect 134 534 270 535
rect 143 526 270 534
rect 295 521 302 523
rect 191 515 302 521
rect 493 483 498 538
rect 552 490 557 553
rect 493 482 508 483
rect 493 478 539 482
rect 109 394 218 400
rect 566 394 571 478
rect 410 389 571 394
rect 120 382 251 383
rect 127 376 251 382
rect 180 367 275 372
rect 299 365 306 366
rect 191 362 195 363
rect 191 358 299 362
rect 191 357 195 358
rect 116 213 201 218
rect 169 194 255 199
rect 177 185 280 190
rect 300 181 308 185
rect 191 174 308 181
rect 127 54 132 58
rect -70 39 -4 42
rect -92 -66 -88 -61
rect -93 -152 -90 -146
rect -84 -231 -81 -226
rect -81 -234 -76 -231
rect -80 -856 -77 -234
rect -70 -372 -67 39
rect 127 -12 131 54
rect 127 -16 230 -12
rect 124 -35 162 -31
rect 168 -35 219 -31
rect -33 -50 -4 -47
rect -33 -61 -30 -50
rect -33 -351 -30 -66
rect 215 -76 219 -35
rect 226 -63 230 -16
rect 226 -67 380 -63
rect 215 -80 224 -76
rect 230 -80 354 -76
rect 376 -78 380 -67
rect 376 -84 378 -78
rect 215 -88 333 -84
rect 126 -125 172 -121
rect 177 -125 194 -121
rect 215 -121 219 -88
rect 200 -125 219 -121
rect 236 -100 298 -96
rect -26 -140 -5 -137
rect -26 -146 -22 -140
rect -26 -336 -22 -152
rect 126 -214 133 -210
rect 236 -210 240 -100
rect 139 -214 242 -210
rect 148 -218 155 -214
rect 134 -222 155 -218
rect -13 -229 -5 -226
rect -26 -340 2 -336
rect -2 -351 2 -340
rect 134 -342 138 -222
rect 192 -339 308 -332
rect 300 -343 308 -339
rect 138 -348 280 -343
rect -33 -353 -25 -351
rect -33 -354 -28 -353
rect 198 -357 255 -352
rect 198 -372 201 -371
rect -70 -375 201 -372
rect 198 -376 201 -375
rect -27 -517 -23 -389
rect -27 -521 -3 -517
rect -7 -538 -3 -521
rect 132 -525 136 -389
rect 204 -520 299 -516
rect 299 -524 306 -523
rect 137 -529 275 -525
rect 196 -530 275 -529
rect 196 -538 251 -534
rect -26 -575 -16 -541
rect -8 -541 251 -538
rect -8 -542 199 -541
rect 410 -552 571 -547
rect 129 -561 137 -554
rect 129 -700 136 -561
rect 566 -636 571 -552
rect 493 -640 539 -636
rect 493 -641 508 -640
rect 205 -679 302 -673
rect 295 -681 302 -679
rect 493 -696 498 -641
rect 129 -707 237 -700
rect 386 -711 391 -710
rect 552 -711 557 -648
rect 386 -715 557 -711
rect 388 -716 557 -715
rect -80 -869 -72 -856
rect 260 -869 265 -866
rect -80 -877 265 -869
rect 493 -878 498 -729
rect 381 -883 498 -878
<< m3contact >>
rect -88 -66 -83 -61
rect -90 -152 -84 -146
rect -81 -231 -76 -226
rect -33 -66 -28 -61
rect -26 -152 -19 -146
rect -18 -231 -13 -226
<< metal3 >>
rect -83 -66 -33 -61
rect -84 -152 -26 -146
rect -76 -231 -18 -226
use XNOR  XNOR_3
timestamp 1701500099
transform 1 0 -13 0 1 -168
box 4 -88 140 -19
use XNOR  XNOR_2
timestamp 1701500099
transform 1 0 -13 0 1 -79
box 4 -88 140 -19
use XNOR  XNOR_1
timestamp 1701500099
transform 1 0 -12 0 1 11
box 4 -88 140 -19
use 4_AND  4_AND_0
timestamp 1700312805
transform 1 0 360 0 1 -65
box -60 -95 126 46
use XNOR  XNOR_0
timestamp 1701500099
transform 1 0 -12 0 1 100
box 4 -88 140 -19
use 5_AND  5_AND_0
timestamp 1699296593
transform 1 0 261 0 1 213
box -60 -99 162 46
use 3_AND  3_AND_0
timestamp 1701512323
transform 1 0 300 0 1 554
box -60 -95 82 46
use 4_AND  4_AND_1
timestamp 1700312805
transform 1 0 280 0 1 391
box -60 -95 126 46
use 4_OR  4_OR_0
timestamp 1699298635
transform 1 0 555 0 1 486
box -44 -48 127 28
use AND  AND_0
timestamp 1700315882
transform 1 0 299 0 1 722
box -60 -96 78 46
<< labels >>
rlabel metal1 -17 -39 -16 -38 3 a1
rlabel metal1 -18 -130 -17 -129 3 a2
rlabel metal1 -18 -218 -17 -217 3 a3
rlabel polycontact 83 -5 84 -4 1 b1_not
rlabel polysilicon 29 -6 30 -5 1 a1_not
rlabel polysilicon 27 -97 28 -96 1 a2_not
rlabel polysilicon 82 -96 83 -95 1 b2_not
rlabel polysilicon 27 -186 28 -185 1 a3_not
rlabel polysilicon 81 -186 82 -185 1 b3_not
rlabel metal1 -17 50 -16 51 3 a0
rlabel metal2 -17 40 -16 41 3 b0
rlabel polysilicon 28 85 29 86 5 a0_not
rlabel polysilicon 83 85 84 86 5 b0_not
rlabel metal1 53 83 54 84 5 vdd
rlabel metal1 53 8 54 10 1 gnd
rlabel metal2 271 -66 274 -64 1 check1
rlabel metal2 269 -79 272 -77 1 check2
rlabel metal2 265 -99 268 -97 1 check4
rlabel metal1 707 472 710 476 7 greater_than
rlabel metal1 604 -66 605 -65 1 equal_to
rlabel metal1 707 -635 710 -633 7 less_than
rlabel metal2 -83 -229 -82 -228 1 b3
rlabel metal2 -92 -150 -91 -148 3 b2
rlabel metal2 -91 -64 -90 -62 3 b1
rlabel metal2 165 -124 169 -122 1 check3
<< end >>
